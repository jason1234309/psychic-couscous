module top(
  input LIOB33_SING_X0Y149_IOB_X0Y149_IPAD,
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_X0Y141_IOB_X0Y141_IPAD,
  input LIOB33_X0Y141_IOB_X0Y142_IPAD,
  input LIOB33_X0Y143_IOB_X0Y143_IPAD,
  input LIOB33_X0Y145_IOB_X0Y145_IPAD,
  input LIOB33_X0Y145_IOB_X0Y146_IPAD,
  input LIOB33_X0Y147_IOB_X0Y147_IPAD,
  input LIOB33_X0Y147_IOB_X0Y148_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y177_IOB_X0Y178_IPAD,
  input LIOB33_X0Y179_IOB_X0Y179_IPAD,
  input LIOB33_X0Y179_IOB_X0Y180_IPAD,
  input LIOB33_X0Y181_IOB_X0Y181_IPAD,
  input LIOB33_X0Y181_IOB_X0Y182_IPAD,
  input LIOB33_X0Y183_IOB_X0Y183_IPAD,
  input LIOB33_X0Y183_IOB_X0Y184_IPAD,
  input LIOB33_X0Y185_IOB_X0Y185_IPAD,
  input LIOB33_X0Y185_IOB_X0Y186_IPAD,
  input LIOB33_X0Y187_IOB_X0Y187_IPAD,
  input LIOB33_X0Y187_IOB_X0Y188_IPAD,
  input LIOB33_X0Y189_IOB_X0Y189_IPAD,
  input LIOB33_X0Y189_IOB_X0Y190_IPAD,
  input LIOB33_X0Y191_IOB_X0Y191_IPAD,
  input LIOB33_X0Y191_IOB_X0Y192_IPAD,
  input LIOB33_X0Y193_IOB_X0Y193_IPAD,
  input LIOB33_X0Y193_IOB_X0Y194_IPAD,
  input LIOB33_X0Y195_IOB_X0Y195_IPAD,
  input LIOB33_X0Y195_IOB_X0Y196_IPAD,
  input LIOB33_X0Y197_IOB_X0Y197_IPAD,
  input LIOB33_X0Y197_IOB_X0Y198_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output RIOB33_SING_X105Y100_IOB_X1Y100_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_X105Y101_IOB_X1Y101_OPAD,
  output RIOB33_X105Y101_IOB_X1Y102_OPAD,
  output RIOB33_X105Y103_IOB_X1Y103_OPAD,
  output RIOB33_X105Y103_IOB_X1Y104_OPAD,
  output RIOB33_X105Y105_IOB_X1Y105_OPAD,
  output RIOB33_X105Y105_IOB_X1Y106_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y113_IOB_X1Y114_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CLK;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_SR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CLK;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_SR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AMUX;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CLK;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CMUX;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_SR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CLK;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_SR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CLK;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_SR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CLK;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_SR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CLK;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_SR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CLK;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_SR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_SR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_SR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_SR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_SR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_SR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_SR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_SR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_SR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_SR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_SR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_SR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_SR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_SR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_SR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_AMUX;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_AO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_AO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_A_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_BO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_B_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_CO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_CO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_C_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_DO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_DO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X12Y100_D_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_AO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_AO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_A_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_BO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_BO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_B_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_CO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_CO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_C_XOR;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D1;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D2;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D3;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D4;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_DO5;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_DO6;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D_CY;
  wire [0:0] CLBLM_L_X10Y100_SLICE_X13Y100_D_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_AMUX;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_AO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_BO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_CO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_DO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_AMUX;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_AO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_BO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_CO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_CO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_DO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_DO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CLK;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_SR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CLK;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_SR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CLK;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_SR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CLK;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_SR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_SR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CLK;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_SR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_SR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_SR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_SR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_SR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_SR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_SR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_SR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_SR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_SR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_SR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_SR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_SR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_SR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_SR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_SR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BMUX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_SR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_SR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_SR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_SR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_SR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_SR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_SR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_SR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_SR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_SR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_SR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_AO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_AO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_A_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_BO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_BO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_B_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_CO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_CO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_C_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_DO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_DO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X16Y100_D_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_AO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_AO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_A_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_BO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_BO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_B_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_CO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_CO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_C_XOR;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D1;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D2;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D3;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D4;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_DO5;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_DO6;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D_CY;
  wire [0:0] CLBLM_L_X12Y100_SLICE_X17Y100_D_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_AMUX;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_AO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_AO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_A_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_BO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_BO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_B_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_CLK;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_CO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_CO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_C_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_DO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_DO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_D_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X16Y101_SR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_AO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_AO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_A_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_BO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_BO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_B_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_CMUX;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_CO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_CO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_C_XOR;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D1;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D2;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D3;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D4;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_DMUX;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_DO5;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_DO6;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D_CY;
  wire [0:0] CLBLM_L_X12Y101_SLICE_X17Y101_D_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_AO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_AO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_A_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_BO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_BO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_B_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_CLK;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_CMUX;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_CO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_CO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_C_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_DO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_DO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_D_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X16Y102_SR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_AMUX;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_AO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_AO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_A_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_BO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_BO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_B_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_CO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_CO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_C_XOR;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D1;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D2;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D3;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D4;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_DO5;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_DO6;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D_CY;
  wire [0:0] CLBLM_L_X12Y102_SLICE_X17Y102_D_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_AO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_AO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_A_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_BMUX;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_BO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_BO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_B_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_CLK;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_CO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_CO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_C_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_DO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_DO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_D_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X16Y103_SR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_AO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_AO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_A_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_BO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_BO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_B_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_CLK;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_CO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_CO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_C_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D1;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D2;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D3;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D4;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_DO5;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_DO6;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D_CY;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_D_XOR;
  wire [0:0] CLBLM_L_X12Y103_SLICE_X17Y103_SR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CLK;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CMUX;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_DO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_SR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_AO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_AO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_BO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_BO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_CO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_CO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_DO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_DO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DMUX;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AMUX;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CLK;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_SR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CLK;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_SR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CLK;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_SR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AMUX;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CLK;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_SR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CLK;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_SR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CLK;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_SR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CLK;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_SR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5Q;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_SR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BMUX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_SR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X16Y116_SR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_A_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_B_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CLK;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CMUX;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_C_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D1;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D2;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D3;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D4;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO5;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_CY;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_D_XOR;
  wire [0:0] CLBLM_L_X12Y116_SLICE_X17Y116_SR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_SR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_SR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_SR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_SR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DMUX;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_SR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X16Y122_SR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_A_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_B_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CLK;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_C_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D1;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D2;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D3;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D4;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DMUX;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO5;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_CY;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_D_XOR;
  wire [0:0] CLBLM_L_X12Y122_SLICE_X17Y122_SR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CMUX;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X16Y123_SR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_A_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_B_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CLK;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_C_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D1;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D2;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D3;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D4;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO5;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_CY;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_D_XOR;
  wire [0:0] CLBLM_L_X12Y123_SLICE_X17Y123_SR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X16Y124_SR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_A_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_B_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CLK;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_C_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D1;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D2;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D3;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D4;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DMUX;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO5;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_CY;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_D_XOR;
  wire [0:0] CLBLM_L_X12Y124_SLICE_X17Y124_SR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CLK;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DMUX;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X16Y125_SR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_A_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_B_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_C_XOR;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D1;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D2;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D3;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D4;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO5;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_CY;
  wire [0:0] CLBLM_L_X12Y125_SLICE_X17Y125_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BMUX;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_SR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_SR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_SR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CMUX;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_SR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_SR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_SR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_SR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_SR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_SR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_SR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_SR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_AO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_AO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_A_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_BMUX;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_BO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_BO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_B_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_CLK;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_CO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_CO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_C_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_DO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_DO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_D_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X22Y101_SR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_AO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_AO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_A_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_BO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_BO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_B_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_CO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_CO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_C_XOR;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D1;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D2;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D3;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D4;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_DO5;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_DO6;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D_CY;
  wire [0:0] CLBLM_L_X16Y101_SLICE_X23Y101_D_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_AO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_AO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_A_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_BMUX;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_BO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_BO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_B_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_CLK;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_CMUX;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_CO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_CO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_C_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_DO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_DO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_D_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X22Y102_SR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_AMUX;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_AO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_AO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_A_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_BO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_BO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_B_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_CO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_CO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_C_XOR;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D1;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D2;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D3;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D4;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_DO5;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_DO6;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D_CY;
  wire [0:0] CLBLM_L_X16Y102_SLICE_X23Y102_D_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_AO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_AO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_A_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_BO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_BO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_B_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_CO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_CO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_C_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_DMUX;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_DO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_DO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X22Y103_D_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_AO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_AO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_A_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_BO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_BO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_B_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_CO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_C_XOR;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D1;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D2;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D3;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D4;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_DO5;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_DO6;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D_CY;
  wire [0:0] CLBLM_L_X16Y103_SLICE_X23Y103_D_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_AO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_AO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_A_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_BO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_BO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_B_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_CLK;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_CO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_CO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_C_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_DO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_DO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_D_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X22Y104_SR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_AO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_AO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_A_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_BO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_BO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_B_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_CLK;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_CO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_CO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_C_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D1;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D2;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D3;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D4;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_DO5;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_DO6;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D_CY;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_D_XOR;
  wire [0:0] CLBLM_L_X16Y104_SLICE_X23Y104_SR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_AO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_AO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_A_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_BO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_BO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_B_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_CLK;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_CO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_CO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_C_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_DO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_DO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_D_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X22Y105_SR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_AMUX;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_AO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_AO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_A_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_BO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_BO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_B_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_CO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_CO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_C_XOR;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D1;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D2;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D3;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D4;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_DO5;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_DO6;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D_CY;
  wire [0:0] CLBLM_L_X16Y105_SLICE_X23Y105_D_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_AO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_AO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_A_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_BMUX;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_BO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_BO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_B_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_CLK;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_CMUX;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_CO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_CO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_C_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_DO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_DO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_D_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X22Y106_SR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_AMUX;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_AO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_AO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_A_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_BMUX;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_BO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_BO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_B_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_CMUX;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_CO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_CO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_C_XOR;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D1;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D2;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D3;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D4;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_DO5;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_DO6;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D_CY;
  wire [0:0] CLBLM_L_X16Y106_SLICE_X23Y106_D_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_AO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_AO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_A_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_BO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_BO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_B_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_CLK;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_CO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_CO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_C_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_DO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_DO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_D_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X22Y107_SR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_AO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_AO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_A_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_BO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_BO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_B_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_CO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_CO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_C_XOR;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D1;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D2;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D3;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D4;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_DMUX;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_DO5;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_DO6;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D_CY;
  wire [0:0] CLBLM_L_X16Y107_SLICE_X23Y107_D_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_AMUX;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_AO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_AO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_A_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_BO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_BO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_B_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_CLK;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_CO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_CO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_C_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_DO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_DO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_D_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X22Y108_SR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_AO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_AO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_A_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_BO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_BO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_B_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_CO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_CO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_C_XOR;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D1;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D2;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D3;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D4;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_DO5;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_DO6;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D_CY;
  wire [0:0] CLBLM_L_X16Y108_SLICE_X23Y108_D_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_AMUX;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_AO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_AO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_A_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_BMUX;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_BO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_BO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_B_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_CO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_CO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_C_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_DO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_DO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X22Y109_D_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_AMUX;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_AO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_AO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_A_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_BO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_BO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_B_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_CO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_CO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_C_XOR;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D1;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D2;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D3;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D4;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_DO5;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_DO6;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D_CY;
  wire [0:0] CLBLM_L_X16Y109_SLICE_X23Y109_D_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_AO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_AO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_A_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_BO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_BO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_B_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_CLK;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_CO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_CO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_C_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_DO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_DO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_D_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X22Y110_SR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_AMUX;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_AO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_A_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_BO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_BO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_B_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_CO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_CO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_C_XOR;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D1;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D2;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D3;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D4;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_DO5;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_DO6;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D_CY;
  wire [0:0] CLBLM_L_X16Y110_SLICE_X23Y110_D_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_AO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_AO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_A_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_BO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_BO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_B_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_CLK;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_CO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_CO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_C_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_DO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_DO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_D_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X22Y111_SR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_AO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_AO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_A_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_BMUX;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_BO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_B_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_CLK;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_CO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_CO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_C_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D1;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D2;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D3;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D4;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_DO5;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_DO6;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D_CY;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_D_XOR;
  wire [0:0] CLBLM_L_X16Y111_SLICE_X23Y111_SR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_AMUX;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_AO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_AO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_A_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_BMUX;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_BO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_BO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_B_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_CMUX;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_CO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_CO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_C_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_DO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_DO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X22Y113_D_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_AO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_AO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_A_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_BO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_BO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_B_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_CO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_CO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_C_XOR;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D1;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D2;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D3;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D4;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_DO5;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_DO6;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D_CY;
  wire [0:0] CLBLM_L_X16Y113_SLICE_X23Y113_D_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_AO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_AO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_AQ;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_A_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_BMUX;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_BO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_BO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_B_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_CLK;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_CMUX;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_CO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_CO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_C_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_DO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_DO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_D_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X22Y114_SR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_AO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_AO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_AQ;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_A_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_BO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_BO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_BQ;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_B_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_CLK;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_CO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_CO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_C_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D1;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D2;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D3;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D4;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_DO5;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_DO6;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D_CY;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_D_XOR;
  wire [0:0] CLBLM_L_X16Y114_SLICE_X23Y114_SR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_AO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_AO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_AQ;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_A_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_BO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_B_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_CLK;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_CO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_CO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_C_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_DO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_DO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_D_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X22Y115_SR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_AO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_AO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_AQ;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_A_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_BO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_BO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_BQ;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_B_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_CLK;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_CMUX;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_CO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_CO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_C_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D1;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D2;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D3;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D4;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_DO5;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_DO6;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D_CY;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_D_XOR;
  wire [0:0] CLBLM_L_X16Y115_SLICE_X23Y115_SR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_AMUX;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_AO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_AO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_A_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_BMUX;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_BO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_BO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_B_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_CMUX;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_CO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_CO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_C_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_DO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_DO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X22Y116_D_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_AO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_AO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_AQ;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_A_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_BO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_BO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_BQ;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_B_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_CLK;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_CO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_CO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_C_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D1;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D2;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D3;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D4;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_DO5;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_DO6;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D_CY;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_D_XOR;
  wire [0:0] CLBLM_L_X16Y116_SLICE_X23Y116_SR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_AO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_AO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_AQ;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_A_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_BO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_BO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_BQ;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_B_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_CLK;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_CO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_CO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_C_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_DO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_DO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_D_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X22Y117_SR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_AMUX;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_AO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_AO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_A_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_BO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_BO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_B_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_CO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_CO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_C_XOR;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D1;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D2;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D3;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D4;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_DO5;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_DO6;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D_CY;
  wire [0:0] CLBLM_L_X16Y117_SLICE_X23Y117_D_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_AO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_AO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_A_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_BO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_BO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_B_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_CO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_CO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_C_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_DO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_DO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X22Y118_D_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_AO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_AO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_A_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_BO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_BO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_B_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_CLK;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_CO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_CO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_C_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D1;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D2;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D3;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D4;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_DO5;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_DO6;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D_CY;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_D_XOR;
  wire [0:0] CLBLM_L_X16Y118_SLICE_X23Y118_SR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_AO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_AO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_AQ;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_A_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_BMUX;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_BO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_BO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_B_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_CLK;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_CMUX;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_CO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_CO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_C_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_DO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_DO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_D_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X22Y119_SR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_AO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_AO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_AQ;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_A_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_BO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_BO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_B_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_CLK;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_CO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_CO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_C_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D1;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D2;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D3;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D4;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_DO5;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_DO6;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D_CY;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_D_XOR;
  wire [0:0] CLBLM_L_X16Y119_SLICE_X23Y119_SR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_AO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_AO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_AQ;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_A_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_BO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_BO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_B_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_CLK;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_CO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_CO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_C_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_DO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_DO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_D_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X22Y121_SR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_AO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_AO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_A_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_BO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_BO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_B_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_CO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_CO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_C_XOR;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D1;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D2;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D3;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D4;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_DO5;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_DO6;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D_CY;
  wire [0:0] CLBLM_L_X16Y121_SLICE_X23Y121_D_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_AMUX;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_AO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_AO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_A_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_BO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_B_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_CO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_CO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_C_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_DO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_DO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X22Y123_D_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_AO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_AO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_A_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_BO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_BO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_B_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_CO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_CO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_C_XOR;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D1;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D2;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D3;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D4;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_DO5;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_DO6;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D_CY;
  wire [0:0] CLBLM_L_X16Y123_SLICE_X23Y123_D_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_AO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_AO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_AQ;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_A_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_BMUX;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_BO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_BO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_B_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_CLK;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_CMUX;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_CO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_CO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_C_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_DO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_D_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X22Y125_SR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_AMUX;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_AO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_AO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_A_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_BO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_B_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_CO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_C_XOR;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D1;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D2;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D3;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D4;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_DO5;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_DO6;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D_CY;
  wire [0:0] CLBLM_L_X16Y125_SLICE_X23Y125_D_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_AO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_AO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_AQ;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_A_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_BMUX;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_BO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_BO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_B_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_CLK;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_CO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_CO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_C_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_DO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_DO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_D_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X22Y126_SR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_AMUX;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_A_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_BMUX;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_B_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_CO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_C_XOR;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D1;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D2;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D3;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D4;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_DO5;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_DO6;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D_CY;
  wire [0:0] CLBLM_L_X16Y126_SLICE_X23Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_AO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_BO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_CO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_DO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AMUX;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_BO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_CO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_DO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CLK;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_SR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CLK;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_SR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BMUX;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CLK;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_SR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CLK;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_SR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CLK;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_SR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CLK;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_SR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CLK;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_SR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CLK;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_SR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CLK;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_SR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_SR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_SR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_SR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_SR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_SR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_SR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_SR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_SR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_SR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AMUX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_SR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_SR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_SR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_SR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_SR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_SR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_SR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_SR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_SR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_SR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_SR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_SR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_SR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_SR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_AMUX;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_AO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_AO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_A_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_BO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_B_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_CO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_CO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_C_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_DO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_DO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X14Y100_D_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_AO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_AO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_A_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_BO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_BO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_B_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_CO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_CO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_C_XOR;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D1;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D2;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D3;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D4;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_DO5;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_DO6;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D_CY;
  wire [0:0] CLBLM_R_X11Y100_SLICE_X15Y100_D_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_AO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_AO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_A_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_BO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_BO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_B_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_CLK;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_CO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_CO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_C_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_DO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_DO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_D_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X14Y101_SR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_AMUX;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_AO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_AO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_A_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_BO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_BO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_B_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_CO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_CO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_C_XOR;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D1;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D2;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D3;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D4;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_DO5;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_DO6;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D_CY;
  wire [0:0] CLBLM_R_X11Y101_SLICE_X15Y101_D_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_AMUX;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_AO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_AO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_A_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_BO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_BO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_B_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_CO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_CO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_C_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_DO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_DO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X14Y102_D_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_AMUX;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_AO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_AO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_A_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_BO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_BO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_B_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_CMUX;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_CO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_CO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_C_XOR;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D1;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D2;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D3;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D4;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_DO5;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_DO6;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D_CY;
  wire [0:0] CLBLM_R_X11Y102_SLICE_X15Y102_D_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_AO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_BO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_BO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_CLK;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_CMUX;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_CO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_CO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_DMUX;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_DO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_SR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_AO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_AO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_BO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_BO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_CO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_CO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_DO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_DO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CLK;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_SR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CLK;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_SR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CLK;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_SR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CLK;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_SR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CLK;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_SR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_SR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_SR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_SR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_SR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_SR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_SR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_SR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_SR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_SR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_SR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_SR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_SR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AMUX;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_SR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_SR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BMUX;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_SR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_SR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_SR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_SR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_SR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_SR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_SR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_SR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_SR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_SR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_SR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_SR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_SR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_AO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_AO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_A_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_BMUX;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_BO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_BO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_B_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_CLK;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_CO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_C_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_DMUX;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_DO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_DO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_D_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X18Y100_SR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_AO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_A_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_BMUX;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_BO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_BO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_B_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_CO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_CO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_C_XOR;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D1;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D2;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D3;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D4;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_DO5;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_DO6;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D_CY;
  wire [0:0] CLBLM_R_X13Y100_SLICE_X19Y100_D_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_AO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_AO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_A_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_BMUX;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_BO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_BO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_B_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_CLK;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_CO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_CO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_C_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_DO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_DO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_D_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X18Y101_SR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_AMUX;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_AO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_AO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_A_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_BO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_BO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_B_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_CO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_CO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_C_XOR;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D1;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D2;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D3;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D4;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_DO5;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D_CY;
  wire [0:0] CLBLM_R_X13Y101_SLICE_X19Y101_D_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_AO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_AO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_A_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_BO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_BO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_B_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_CLK;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_CMUX;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_CO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_CO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_C_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_DO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_DO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_D_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X18Y102_SR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_AMUX;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_AO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_AO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_A_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_BO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_BO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_B_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_CO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_CO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_C_XOR;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D1;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D2;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D3;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D4;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_DO5;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_DO6;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D_CY;
  wire [0:0] CLBLM_R_X13Y102_SLICE_X19Y102_D_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_AO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_AO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_A_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_BMUX;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_BO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_BO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_B_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_CLK;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_CO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_CO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_C_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_DO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_DO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_D_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X18Y103_SR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_AMUX;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_AO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_AO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_A_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_BO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_BO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_B_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_CO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_CO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_C_XOR;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D1;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D2;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D3;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D4;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_DO5;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_DO6;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D_CY;
  wire [0:0] CLBLM_R_X13Y103_SLICE_X19Y103_D_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_AO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_AO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_A_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_BO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_BO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_B_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_CLK;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_CO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_CO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_C_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_DO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_DO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_D_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X18Y104_SR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_AO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_AO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_A_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_BO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_BO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_B_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_CLK;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_CO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_CO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_C_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D1;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D2;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D3;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D4;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_DO5;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_DO6;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D_CY;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_D_XOR;
  wire [0:0] CLBLM_R_X13Y104_SLICE_X19Y104_SR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AMUX;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_BO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_CO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_DO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_DO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_DO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AMUX;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_DO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_DO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CLK;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_SR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AMUX;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DMUX;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CLK;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_SR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_A_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BMUX;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_B_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CLK;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_C_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DMUX;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X18Y111_SR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_A_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_B_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_C_XOR;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D1;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D2;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D3;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D4;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_DO5;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_DO6;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D_CY;
  wire [0:0] CLBLM_R_X13Y111_SLICE_X19Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CLK;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_SR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AMUX;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CLK;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_SR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_AMUX;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_AO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_AO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_A_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_BO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_BO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_B_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_CO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_CO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_C_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_DO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_DO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X18Y114_D_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_AMUX;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_AO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_AO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_A_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_BO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_B_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_CLK;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_CO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_CO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_C_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D1;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D2;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D3;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D4;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_DO5;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_DO6;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D_CY;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_D_XOR;
  wire [0:0] CLBLM_R_X13Y114_SLICE_X19Y114_SR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AMUX;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_A_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_B_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CLK;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_C_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_DO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_D_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X18Y115_SR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_A_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_BO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_B_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_C_XOR;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D1;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D2;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D3;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D4;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_DO5;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D_CY;
  wire [0:0] CLBLM_R_X13Y115_SLICE_X19Y115_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CLK;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_SR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AMUX;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BMUX;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CLK;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_DO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_SR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_DO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_DO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CLK;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_SR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CLK;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CMUX;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_SR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CLK;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X18Y121_SR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_A_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_B_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CLK;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_C_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D1;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D2;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D3;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D4;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO5;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_CY;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_D_XOR;
  wire [0:0] CLBLM_R_X13Y121_SLICE_X19Y121_SR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X18Y122_SR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_A_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_B_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CLK;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_C_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D1;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D2;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D3;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D4;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO5;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_CY;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_D_XOR;
  wire [0:0] CLBLM_R_X13Y122_SLICE_X19Y122_SR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X18Y123_SR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_A_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_B_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CLK;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_C_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D1;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D2;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D3;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D4;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO5;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_CY;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_D_XOR;
  wire [0:0] CLBLM_R_X13Y123_SLICE_X19Y123_SR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_BQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CLK;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X18Y124_SR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_A_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BMUX;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_B_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CLK;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_C_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D1;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D2;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D3;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D4;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO5;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_CY;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_D_XOR;
  wire [0:0] CLBLM_R_X13Y124_SLICE_X19Y124_SR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BMUX;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X18Y125_SR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_A_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_B_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CLK;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_C_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D1;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D2;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D3;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D4;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO5;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_CY;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_D_XOR;
  wire [0:0] CLBLM_R_X13Y125_SLICE_X19Y125_SR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X18Y126_SR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_A_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_B_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CLK;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_C_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D1;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D2;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D3;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D4;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO5;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_CY;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_D_XOR;
  wire [0:0] CLBLM_R_X13Y126_SLICE_X19Y126_SR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CLK;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_SR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CLK;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_SR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CLK;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_SR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_SR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_SR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_SR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BMUX;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_SR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CLK;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_SR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AMUX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_AO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_AO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_A_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_BMUX;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_BO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_BO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_B_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_CLK;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_CO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_CO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_C_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_DMUX;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_DO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_DO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_D_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X20Y100_SR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_AO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_AO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_A_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_BO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_BO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_B_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_CO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_C_XOR;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D1;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D2;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D3;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D4;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_DO5;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_DO6;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D_CY;
  wire [0:0] CLBLM_R_X15Y100_SLICE_X21Y100_D_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_AMUX;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_AO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_A_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_BMUX;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_BO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_BO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_B_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_CO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_CO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_C_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_DO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_DO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X20Y101_D_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_AMUX;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_AO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_AO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_A_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_BMUX;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_BO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_BO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_B_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_CO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_CO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_C_XOR;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D1;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D2;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D3;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D4;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_DO5;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_DO6;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D_CY;
  wire [0:0] CLBLM_R_X15Y101_SLICE_X21Y101_D_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_AO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_AO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_A_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_BO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_BO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_B_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_CLK;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_CO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_CO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_C_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_DO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_DO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_D_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X20Y102_SR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_AMUX;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_AO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_AO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_A_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_BO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_B_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_CO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_CO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_C_XOR;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D1;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D2;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D3;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D4;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_DO5;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_DO6;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D_CY;
  wire [0:0] CLBLM_R_X15Y102_SLICE_X21Y102_D_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_AMUX;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_AO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_AO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_A_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_BO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_BO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_B_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_CMUX;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_CO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_CO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_C_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_DO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_DO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X20Y103_D_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_AMUX;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_AO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_AO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_A_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_BO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_BO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_B_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_CO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_CO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_C_XOR;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D1;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D2;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D3;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D4;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_DO5;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_DO6;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D_CY;
  wire [0:0] CLBLM_R_X15Y103_SLICE_X21Y103_D_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_AO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_AO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_A_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_BO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_BO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_B_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_CLK;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_CO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_CO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_C_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_DO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_DO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_D_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X20Y104_SR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_AO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_AO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_A_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_BO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_BO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_B_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_CLK;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_CO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_CO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_C_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D1;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D2;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D3;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D4;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_DO5;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_DO6;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D_CY;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_D_XOR;
  wire [0:0] CLBLM_R_X15Y104_SLICE_X21Y104_SR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_AO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_AO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_A_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_BO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_BO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_B_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_CO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_CO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_C_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_DMUX;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_DO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_DO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X20Y105_D_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_AO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_AO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_A_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_BMUX;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_BO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_BO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_B_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_CLK;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_CO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_CO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_C_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D1;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D2;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D3;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D4;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_DO5;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_DO6;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D_CY;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_D_XOR;
  wire [0:0] CLBLM_R_X15Y105_SLICE_X21Y105_SR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_AO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_AO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_A_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_BO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_BO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_B_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_CLK;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_CO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_CO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_C_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_DMUX;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_DO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_DO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_D_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X20Y106_SR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_AO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_AO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_A_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_BMUX;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_BO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_BO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_B_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_CO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_CO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_C_XOR;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D1;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D2;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D3;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D4;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_DO5;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_DO6;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D_CY;
  wire [0:0] CLBLM_R_X15Y106_SLICE_X21Y106_D_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_AO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_AO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_A_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_BMUX;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_BO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_BO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_B_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_CLK;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_CMUX;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_CO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_CO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_C_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_DO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_DO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_D_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X20Y107_SR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_AMUX;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_AO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_AO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_A_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_BO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_BO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_B_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_CLK;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_CO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_CO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_CQ;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_C_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D1;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D2;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D3;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D4;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_DO5;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_DO6;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D_CY;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_D_XOR;
  wire [0:0] CLBLM_R_X15Y107_SLICE_X21Y107_SR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_AMUX;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_AO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_AO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_A_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_BO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_BO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_B_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_CO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_CO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_C_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_DO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_DO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X20Y108_D_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_AMUX;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_AO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_AO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_A_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_BO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_BO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_B_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_CO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_CO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_C_XOR;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D1;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D2;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D3;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D4;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_DMUX;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_DO5;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_DO6;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D_CY;
  wire [0:0] CLBLM_R_X15Y108_SLICE_X21Y108_D_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_AO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_A_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_BO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_B_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_CMUX;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_CO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_CO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_C_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_DO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_DO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X20Y109_D_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_AMUX;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_AO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_AO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_A_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_BO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_BO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_B_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_CO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_CO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_C_XOR;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D1;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D2;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D3;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D4;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_DO5;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_DO6;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D_CY;
  wire [0:0] CLBLM_R_X15Y109_SLICE_X21Y109_D_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_AMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_AO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_A_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_BO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_B_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_CO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_C_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_DO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X20Y110_D_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_AMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_AO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_A_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_BMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_BO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_B_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_CMUX;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_CO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_C_XOR;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D1;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D2;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D3;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D4;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_DO5;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D_CY;
  wire [0:0] CLBLM_R_X15Y110_SLICE_X21Y110_D_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_AMUX;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_AO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_AO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_A_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_BO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_B_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_CO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_CO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_C_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_DMUX;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_DO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_DO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X20Y111_D_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_AO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_AO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_A_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_BO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_B_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_CLK;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_CO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_CO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_C_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D1;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D2;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D3;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D4;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_DO5;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_DO6;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D_CY;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_D_XOR;
  wire [0:0] CLBLM_R_X15Y111_SLICE_X21Y111_SR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_AMUX;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_AO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_AO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_A_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_BO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_BO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_B_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_CO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_CO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_C_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_DO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_DO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X20Y112_D_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_AO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_AO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_A_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_BMUX;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_BO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_B_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_CLK;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_CMUX;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_CO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_CO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_C_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D1;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D2;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D3;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D4;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_DO5;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_DO6;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D_CY;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_D_XOR;
  wire [0:0] CLBLM_R_X15Y112_SLICE_X21Y112_SR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_AO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_A_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_BO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_BO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_B_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_CO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_C_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_DO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X20Y113_D_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_AO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_A_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_BO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_B_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_CO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_C_XOR;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D1;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D2;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D3;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D4;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_DO5;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D_CY;
  wire [0:0] CLBLM_R_X15Y113_SLICE_X21Y113_D_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_AO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_AO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_AQ;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_A_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_BMUX;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_BO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_B_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_CLK;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_CO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_C_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_DO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_D_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X20Y114_SR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_AO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_AO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_AQ;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_A_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_BMUX;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_BO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_BO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_B_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_CLK;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_CO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_C_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D1;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D2;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D3;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D4;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_DO5;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_DO6;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D_CY;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_D_XOR;
  wire [0:0] CLBLM_R_X15Y114_SLICE_X21Y114_SR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_AO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_AO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_AQ;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_A_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_BMUX;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_BO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_BO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_B_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_CLK;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_CO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_CO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_C_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_DO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_DO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_D_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X20Y115_SR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_AO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_AO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_AQ;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_A_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_BO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_BO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_B_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_CLK;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_CMUX;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_CO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_CO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_C_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D1;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D2;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D3;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D4;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_DO5;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D_CY;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_D_XOR;
  wire [0:0] CLBLM_R_X15Y115_SLICE_X21Y115_SR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_AO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_AO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_AQ;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_A_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_BO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_BO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_BQ;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_B_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_CLK;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_CMUX;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_CO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_CO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_C_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_DO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_DO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_D_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X20Y116_SR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_AO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_AO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_AQ;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_A_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_BO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_BO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_BQ;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_B_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_CLK;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_CO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_CO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_C_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D1;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D2;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D3;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D4;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_DO5;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_DO6;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D_CY;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_D_XOR;
  wire [0:0] CLBLM_R_X15Y116_SLICE_X21Y116_SR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_AO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_AO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_AQ;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_A_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_BMUX;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_BO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_BO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_B_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_CLK;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_CMUX;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_CO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_CO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_C_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_DO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_DO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_D_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X20Y117_SR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_AO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_AO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_AQ;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_A_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_BO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_BO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_BQ;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_B_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_CLK;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_CO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_CO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_C_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D1;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D2;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D3;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D4;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_DO5;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_DO6;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D_CY;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_D_XOR;
  wire [0:0] CLBLM_R_X15Y117_SLICE_X21Y117_SR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_AO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_AO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_AQ;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_A_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_BMUX;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_BO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_BO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_B_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_CLK;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_CO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_CO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_C_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_DO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_DO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_D_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X20Y118_SR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_AO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_AO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_AQ;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_A_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_BO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_BO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_B_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_CLK;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_CO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_CO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_C_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D1;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D2;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D3;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D4;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_DO5;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_DO6;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D_CY;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_D_XOR;
  wire [0:0] CLBLM_R_X15Y118_SLICE_X21Y118_SR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_AO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_AO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_AQ;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_A_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_BMUX;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_BO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_BO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_B_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_CLK;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_CMUX;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_CO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_CO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_C_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_DO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_DO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_D_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X20Y119_SR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_AO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_AO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_AQ;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_A_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_BO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_BO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_BQ;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_B_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_CLK;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_CMUX;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_CO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_CO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_C_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D1;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D2;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D3;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D4;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_DO5;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_DO6;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D_CY;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_D_XOR;
  wire [0:0] CLBLM_R_X15Y119_SLICE_X21Y119_SR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_AO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_AO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_AQ;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_A_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_BO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_BO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_B_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_CLK;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_CO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_CO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_C_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_DO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_DO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_D_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X20Y120_SR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_AO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_AO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_AQ;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_A_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_BMUX;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_BO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_B_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_CLK;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_CO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_CO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_C_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D1;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D2;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D3;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D4;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_DO5;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_DO6;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D_CY;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_D_XOR;
  wire [0:0] CLBLM_R_X15Y120_SLICE_X21Y120_SR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_AO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_AO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_AQ;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_A_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_BO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_BO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_BQ;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_B_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_CLK;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_CO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_CO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_C_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_DO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_DO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_D_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X20Y121_SR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_AO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_AO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_AQ;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_A_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_BO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_BO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_B_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_CLK;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_CO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_CO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_C_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D1;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D2;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D3;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D4;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_DO5;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_DO6;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D_CY;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_D_XOR;
  wire [0:0] CLBLM_R_X15Y121_SLICE_X21Y121_SR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_AO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_AQ;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_A_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_BO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_BO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_BQ;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_B_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_CLK;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_CMUX;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_CO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_CO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_C_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_DMUX;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_DO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_DO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_D_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X20Y122_SR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_AO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_AO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_AQ;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_A_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_BO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_BO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_B_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_CLK;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_CO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_CO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_C_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D1;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D2;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D3;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D4;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_DO5;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_DO6;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D_CY;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_D_XOR;
  wire [0:0] CLBLM_R_X15Y122_SLICE_X21Y122_SR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_AO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_AQ;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_A_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_BMUX;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_BO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_BO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_B_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_CLK;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_CMUX;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_CO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_CO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_C_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_DO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_DO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_D_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X20Y123_SR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_AO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_AO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_AQ;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_A_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_BMUX;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_BO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_BO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_B_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_CLK;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_CMUX;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_CO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_CO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_C_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D1;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D2;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D3;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D4;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_DO5;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_DO6;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D_CY;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_D_XOR;
  wire [0:0] CLBLM_R_X15Y123_SLICE_X21Y123_SR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_AO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_AO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_AQ;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_A_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_BMUX;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_BO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_BO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_B_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_CLK;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_CMUX;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_CO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_CO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_C_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_DO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_DO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_D_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X20Y124_SR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_AO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_AO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_AQ;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_A_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_BO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_BO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_B_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_CLK;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_CO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_CO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_C_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D1;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D2;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D3;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D4;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_DO5;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_DO6;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D_CY;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_D_XOR;
  wire [0:0] CLBLM_R_X15Y124_SLICE_X21Y124_SR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_AO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_AO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_A_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_BO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_BO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_B_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_CO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_CO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_C_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_DO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_DO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X20Y125_D_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_AO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_AO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_AQ;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_A_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_BO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_BO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_BQ;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_B_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_CLK;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_CMUX;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_CO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_CO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_C_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D1;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D2;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D3;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D4;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_DO5;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_DO6;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D_CY;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_D_XOR;
  wire [0:0] CLBLM_R_X15Y125_SLICE_X21Y125_SR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_AO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_AO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_AQ;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_A_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_BO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_BO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_BQ;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_B_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_CLK;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_CO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_CO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_C_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_DO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_DO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_D_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X20Y126_SR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_AO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_AO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_AQ;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_A_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_BO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_BO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_B_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_CLK;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_CO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_CO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_C_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D1;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D2;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D3;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D4;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_DMUX;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_DO5;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D_CY;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_D_XOR;
  wire [0:0] CLBLM_R_X15Y126_SLICE_X21Y126_SR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_AO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_AO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_AQ;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_A_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_BO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_BO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_B_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_CLK;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_CO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_CO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_C_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_DO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_DO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_D_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X20Y127_SR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_AMUX;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_AO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_AO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_A_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_BO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_B_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_CO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_C_XOR;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D1;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D2;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D3;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D4;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_DO5;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D_CY;
  wire [0:0] CLBLM_R_X15Y127_SLICE_X21Y127_D_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AMUX;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BMUX;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_DO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AMUX;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_BO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_CO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_DO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CLK;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_DO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_SR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AMUX;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CMUX;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_DO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CLK;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_DO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_SR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CLK;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_DO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_SR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CLK;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_DMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_DO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_DO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_SR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_BO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_BQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CLK;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_DO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_DO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_SR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_AO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_AO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_A_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_BO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_BO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_B_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_CO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_CO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_C_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_DO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_DO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X20Y132_D_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_AO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_AO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_AQ;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_A_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_BO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_BO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_BQ;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_B_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_CLK;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_CO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_CO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_CQ;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_C_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D1;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D2;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D3;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D4;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_DO5;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_DO6;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_DQ;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D_CY;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_D_XOR;
  wire [0:0] CLBLM_R_X15Y132_SLICE_X21Y132_SR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_SR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_SR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_SR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_SR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_SR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_SR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_SR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_SR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_SR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_SR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_SR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_SR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_SR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_SR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_SR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_SR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_SR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_SR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_SR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_SR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_SR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_SR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_SR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CLK;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_SR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CLK;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_SR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CLK;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_SR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_SR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_SR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_SR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CLK;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_SR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_SR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_SR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_SR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_SR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_SR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_SR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_SR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_SR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_SR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_SR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_SR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_SR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_SR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_SR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_SR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_SR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_SR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_I;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_D;
  wire [0:0] LIOI3_SING_X0Y149_ILOGIC_X0Y149_O;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y148_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_O;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccfcccfa0afa0a)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_BQ),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefececa3a3a0a0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_B5Q),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_DO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_BQ),
.I2(CLBLL_L_X2Y116_SLICE_X0Y116_A5Q),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_A5Q),
.I1(CLBLL_L_X2Y116_SLICE_X0Y116_BO6),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedcfedcba10ba10)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.Q(CLBLL_L_X2Y116_SLICE_X0Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.Q(CLBLL_L_X2Y116_SLICE_X0Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecafecafeca0eca0)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y116_SLICE_X0Y116_AQ),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf88b88fbf88b88)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I3(CLBLL_L_X2Y116_SLICE_X0Y116_A5Q),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeccff55eeccaa00)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(CLBLL_L_X2Y116_SLICE_X0Y116_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLL_L_X2Y116_SLICE_X0Y116_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I4(CLBLL_L_X2Y116_SLICE_X0Y116_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.Q(CLBLL_L_X2Y117_SLICE_X0Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffba30ffffba30)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff00aa80ffc0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.Q(CLBLL_L_X2Y117_SLICE_X1Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000077077707)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55055505dd0d5505)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I4(LIOB33_X0Y159_IOB_X0Y160_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.Q(CLBLL_L_X2Y118_SLICE_X0Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y118_SLICE_X0Y118_BO6),
.Q(CLBLL_L_X2Y118_SLICE_X0Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdcdcffff5050)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcceecceeccee)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0a0a0a0bbaaaaaa)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd0ddd0ddd0ddd0d)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.Q(CLBLL_L_X2Y118_SLICE_X1Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeaea0000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f4f0000bfff)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_DO6),
.I5(LIOB33_X0Y151_IOB_X0Y151_I),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a0a0a0a0a0a0a0)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfc0cfca)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y153_I),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.Q(CLBLL_L_X2Y119_SLICE_X0Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd0000d000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(LIOB33_X0Y193_IOB_X0Y194_I),
.I2(LIOB33_X0Y153_IOB_X0Y153_I),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c80cc00dfecffcc)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc33cc33cc3)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0f0000ff0f)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3ffc30000ffc3)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaff0a0fffff0f0f)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696696996966969)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffff70807788)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h11f122f222f222f2)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee0f0effff0f0f)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0aff0aff0a)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h135733ff20aa0000)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ffaa)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff33cc)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I2(1'b1),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000066996996)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1bb212227bbb1bb2)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500ff55f6e2e260)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffacffaca0aca0ac)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8bbf8bbf888f888)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_A5Q),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f5a0f5a0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0f0aaaaf3f0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00eeee)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444fefe5454)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3b3b3b3a0a0a0a0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfc55005d0c5500)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.I1(LIOB33_X0Y161_IOB_X0Y161_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33f030ff33fa32)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(LIOB33_X0Y161_IOB_X0Y161_I),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf033fc33)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(LIOB33_X0Y141_IOB_X0Y141_I),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfcccffcccccc)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000003fffff)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ff4044f0ff)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000051f351f3)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefff0f0f44000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I3(LIOB33_X0Y185_IOB_X0Y185_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(LIOB33_X0Y155_IOB_X0Y155_I),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha088a088ffffa088)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(LIOB33_X0Y159_IOB_X0Y159_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7707550555055505)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I4(LIOB33_X0Y163_IOB_X0Y163_I),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb33bb00aa00aa)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(LIOB33_X0Y161_IOB_X0Y162_I),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555515555555)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555df7ff00000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I4(LIOB33_X0Y161_IOB_X0Y162_I),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaff22332233)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8f0f0fdd880000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I3(LIOB33_X0Y155_IOB_X0Y156_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000080000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa3232fffa3332)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I3(LIOB33_X0Y155_IOB_X0Y156_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc00fcfefe00fe)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(LIOB33_X0Y159_IOB_X0Y159_I),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f21122f1f21122)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc50dca0ec00cc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I5(LIOB33_X0Y157_IOB_X0Y157_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00be3cfaf0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffa2f3a0f0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfceccceccc)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000001f3f1f3f)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fff30ff0fff00)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I5(LIOB33_X0Y163_IOB_X0Y164_I),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c0faf0ccccffff)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ffff0000ffff000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff8f00000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf0000af00)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y146_I),
.I1(1'b1),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_X0Y181_IOB_X0Y181_I),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heecc0e0ceecc0e0c)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(LIOB33_X0Y161_IOB_X0Y161_I),
.I2(LIOB33_X0Y161_IOB_X0Y162_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y159_IOB_X0Y160_I),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffe)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(LIOB33_X0Y159_IOB_X0Y159_I),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(LIOB33_X0Y157_IOB_X0Y158_I),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_DO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_CO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_BO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_AO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_DO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I2(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_CO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55557fd500003fc0)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I5(CLBLM_L_X8Y101_SLICE_X11Y101_CO6),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_BO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880066aa66aa)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_AO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.Q(CLBLM_L_X8Y102_SLICE_X10Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I1(CLBLM_L_X8Y101_SLICE_X11Y101_AO5),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I5(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800080000000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_CLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000080000000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5f5f5a0)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I5(CLBLM_L_X8Y103_SLICE_X11Y103_CO6),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.Q(CLBLM_L_X8Y102_SLICE_X11Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d0c5d0c5d0c5d0c)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_L_X8Y101_SLICE_X11Y101_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1122ffff11221122)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_BLUT (
.I0(CLBLM_L_X10Y101_SLICE_X13Y101_AO5),
.I1(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.I2(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.I4(CLBLM_L_X8Y101_SLICE_X11Y101_CO6),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe3332fffe3332)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y101_SLICE_X11Y101_BO6),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.Q(CLBLM_L_X8Y103_SLICE_X10Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0f33003f0f3300)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00660066ffff0066)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h221111220ff00ff0)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55ff55ee44)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.I2(1'b1),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.Q(CLBLM_L_X8Y103_SLICE_X11Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_DLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff8fff88)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_DO6),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff22fff2)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X11Y103_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5a0f5e4)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I3(CLBLM_L_X8Y103_SLICE_X11Y103_BO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffaafff0ff00)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I1(1'b1),
.I2(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h337b337b005a005a)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf40fd02eaaaaaa8)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I4(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff037503750)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I2(CLBLM_R_X7Y105_SLICE_X9Y105_DO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1177ee88ffff0000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h566aaaaaaaaaaaaa)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa6aaa6aaaaaaa)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_DO6),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h556666aa5a7878f0)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088ccaaff)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccc80000000)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bd004200960096)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800078f078f0)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.Q(CLBLM_L_X8Y105_SLICE_X11Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff00fffcffcc)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_CO6),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f531f531)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fcfcf0000cccc)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555111100550011)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y105_SLICE_X9Y105_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1e875a0f781ef05a)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf531f500f5f5f5f5)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.Q(CLBLM_L_X8Y106_SLICE_X11Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ccfc4454)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfeffffccee)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3f0fffffbfa)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff0fff044)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffc00fd00fc)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050000)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeefeaafa)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff75ff30)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f5500af0faa00)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00aaf0fa)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeff0cffeaffc0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbbbfbbafaaafaa)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0f0f4)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcfeeccfefceecc)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaaae)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff5fff5fff5fff)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5f5fffff5f5f)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0f5f0f1f0f5)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3077f0ffc0c80000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fff7fff7fff7ff)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000000c)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00000066cccccc)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0054ffff4444)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0100ffff0000)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(LIOB33_X0Y185_IOB_X0Y185_I),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1f0a0b1b5a0a0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5530103010)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdffff)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aa00000010)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaafaaaaaaab)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aa000000aa00000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0c0c0c0eac0c0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I5(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0fbfaf3300bbaa)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeafbea51405140)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I4(1'b1),
.I5(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X11Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffae0ceac0)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500330f0efaca)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0fff0aaf000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44440000ff44ff00)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I1(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0cf848fc0cf0c0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000d75f5f5f)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fffff00e2e2)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e4e4e4effffffff)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeccccccfeccfe)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haffacffaaccacaca)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeddeeddcccccccc)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf050f050fff5fff5)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8844221111228844)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa88aa00aa8a)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4fdfdfdf4fdf4)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffaf25af05a)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffafefefafa)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I1(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fffff7f3ffff)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.I2(CLBLM_R_X13Y112_SLICE_X18Y112_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33ff333733)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055ff5557)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000001000)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f800880000)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeef)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(LIOB33_X0Y185_IOB_X0Y185_I),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfcbddcbcfcbcdcb)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(LIOB33_X0Y185_IOB_X0Y185_I),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb8bbbb88b8bbbb)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff50aafa0050)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_DO6),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff404ff0ff404)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_A5Q),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00fff0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f0f0f0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfffffffdff)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h050f050f050f0103)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff222f222)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cc4ecc5f)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdc00dcffdc00dc)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000330033)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I2(1'b1),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafafafaf)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f8f8bbbb8888)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000101fffffefe)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdecfdecb1a0b1a0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fff4f4f4f4f4)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaaeeaa00000000)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_DO6),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.I4(LIOB33_X0Y185_IOB_X0Y185_I),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22fe32ee22fe32)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeaaeeeeaaaa)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf400f000f4f4f0f0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffff88a8ccfc)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.I2(LIOB33_X0Y165_IOB_X0Y166_I),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999988778877)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dddddd00dddddd)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(LIOB33_X0Y151_IOB_X0Y151_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(1'b1),
.I3(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3a3a0000c5c500ff)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaa00aa00aa00)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(LIOB33_X0Y157_IOB_X0Y157_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555505555555)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c0c0c0c0c0c0c0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa0f0afffe0f0e)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I1(LIOB33_X0Y173_IOB_X0Y173_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbaaaa33330000)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(LIOB33_X0Y155_IOB_X0Y156_I),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y171_IOB_X0Y172_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222ff22ff22)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(LIOB33_X0Y175_IOB_X0Y175_I),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0037003f003f003f)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbff0b0faaff0a0f)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22ff222222ff2222)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.I2(1'b1),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(LIOB33_X0Y173_IOB_X0Y174_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0105555505055555)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcffdcff0000dcff)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0ffffa0a0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(LIOB33_X0Y151_IOB_X0Y151_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y167_IOB_X0Y167_I),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ccccff00cc33)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffc0eaf3fb)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(LIOB33_X0Y151_IOB_X0Y152_I),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ffbb5511)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11bb11ffffbb11)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3eef322c0eec022)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111bbbb05af05af)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0f0eeff)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff0fcaaee)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffaa55115500)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I5(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0350035ff350f35f)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h550f3300550f33ff)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000eefeeefe)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_BO6),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_DO6),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff444f4)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I5(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffc0f000f0c)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaaaacfcfcccc)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I3(1'b1),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbf3eac0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I1(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_CO6),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff50f05fff00f00)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I5(LIOB33_X0Y155_IOB_X0Y156_I),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000ddd0d)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(LIOB33_X0Y155_IOB_X0Y155_I),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f044fff0f044ff)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X10Y128_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcba30fcfc3030)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0eac0c0f3fbf3f3)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I2(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafa3afa0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y188_I),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfa0f0f0b0a)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_DO6),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_AO6),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000008caf0405)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I2(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_CO6),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00ff0fff)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000800fffffeff)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X11Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000400fffffffe)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacacacfcacf)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f53705)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I2(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffaffbbbfaaa)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I2(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0fccafee)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(LIOB33_X0Y153_IOB_X0Y153_I),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff737fffff505)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I2(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafa0afa0a0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfe0efc0cfe0e)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y100_SLICE_X12Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y100_SLICE_X12Y100_DO5),
.O6(CLBLM_L_X10Y100_SLICE_X12Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03300330ffff0330)
  ) CLBLM_L_X10Y100_SLICE_X12Y100_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_L_X10Y100_SLICE_X12Y100_AO5),
.I4(CLBLM_L_X10Y101_SLICE_X13Y101_AO5),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_L_X10Y100_SLICE_X12Y100_CO5),
.O6(CLBLM_L_X10Y100_SLICE_X12Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y100_SLICE_X12Y100_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I4(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.O5(CLBLM_L_X10Y100_SLICE_X12Y100_BO5),
.O6(CLBLM_L_X10Y100_SLICE_X12Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c000c000)
  ) CLBLM_L_X10Y100_SLICE_X12Y100_ALUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y100_SLICE_X12Y100_AO5),
.O6(CLBLM_L_X10Y100_SLICE_X12Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y100_SLICE_X13Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y100_SLICE_X13Y100_DO5),
.O6(CLBLM_L_X10Y100_SLICE_X13Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y100_SLICE_X13Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y100_SLICE_X13Y100_CO5),
.O6(CLBLM_L_X10Y100_SLICE_X13Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y100_SLICE_X13Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y100_SLICE_X13Y100_BO5),
.O6(CLBLM_L_X10Y100_SLICE_X13Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y100_SLICE_X13Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y100_SLICE_X13Y100_AO5),
.O6(CLBLM_L_X10Y100_SLICE_X13Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h222f222f2f222f22)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_DLUT (
.I0(CLBLM_R_X11Y100_SLICE_X14Y100_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I3(CLBLM_L_X10Y101_SLICE_X12Y101_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_DO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000080000000)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_CLUT (
.I0(CLBLM_L_X8Y101_SLICE_X11Y101_AO6),
.I1(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_BO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_CO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2800000000000000)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_BLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I2(CLBLM_L_X10Y100_SLICE_X12Y100_AO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_BO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I1(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_AO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_DO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_CO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_BO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h808080806c6c6c6c)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_ALUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_AO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.Q(CLBLM_L_X10Y102_SLICE_X12Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500ffff55005500)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I5(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0880000000000000)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I2(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I5(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffe33323332)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I3(CLBLM_L_X10Y100_SLICE_X12Y100_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000066cccccc)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800800000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I1(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I4(CLBLM_L_X10Y102_SLICE_X13Y102_DO6),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I4(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a00000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.Q(CLBLM_L_X10Y103_SLICE_X12Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f4f4f4f44444444)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_AO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc6ccc6ccccccc)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_CLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_CO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h13ecff007f80ff00)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe00fefffe00fe)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_ALUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_DO6),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I5(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000800000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I1(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_CO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaaaaaaaaaaaaa8)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I5(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccc80000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.Q(CLBLM_L_X10Y104_SLICE_X12Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffa0ffec)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafefefffafffe)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b0d040209060906)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffba5510)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I2(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.Q(CLBLM_L_X10Y104_SLICE_X13Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafefafffffefa)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_DLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2122222222222212)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccfcffffeefe)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_BLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffba5510)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I2(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000000aa000000)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5050ffffdcdc)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ffeaffeaffc0)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7530ba307530ba30)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5ade00cc)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I2(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bb33bb30aa00aa0)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000000)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I1(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000010)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h60ff606088888888)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777888888000000)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccccc)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0f0f2)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333000055005500)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffceffffff0a)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff75ff03)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f066aaaaaa)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff2ffffff22)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff222277a7)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff0080000000)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffce0a)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000010)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffeeffeeeeefef)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I2(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I3(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80010000c0030000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb22ee22ee22ee)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I2(1'b1),
.I3(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff2ffffff22)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafaaefbb)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a0000000800000)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff8fff8f8)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaaa82008282)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaeabeeef)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I2(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff335511ff335511)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfeffffccee)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777752222222)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc5ade00ccf0fc)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4404000044404440)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I3(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h303030ff303030ff)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f01000e0f)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000101111101110)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I2(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I4(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4fff4ff0000f4ff)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000c400c4)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2aaaaaaa80000000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habafaeaa030f0c00)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc00440044)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c5dc0d55d0cd5c0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffaafeab)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff0a0feeff0e0f)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af05af0f0f0f0f0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000010020000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3bffffff0a0a)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffba5510fffa5550)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddddffddff)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.I2(1'b1),
.I3(LIOB33_X0Y185_IOB_X0Y185_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeffffffeedd)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22ff22222fff2f2f)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcff1033cdff0133)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_BO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f441f44ffff1f44)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h75757ff530303ff0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffffc00fcfc)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccdcdccdcf)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f500f5f5f531)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.I4(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_DO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff3f3030f0303)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_CO6),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f0f0fffff0ff)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcfc1030fefe3232)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00010000fffeeebb)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf8fcf8fcf)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(LIOB33_X0Y185_IOB_X0Y185_I),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1fff1fffffffffff)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(LIOB33_X0Y185_IOB_X0Y185_I),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff575555ffff5555)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I2(LIOB33_X0Y185_IOB_X0Y185_I),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff01ff00ff02)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I4(LIOB33_X0Y185_IOB_X0Y185_I),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80808080c0c0f0f0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.I5(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he6f7ccccc0f3cccc)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I5(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfcdcdc)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h303030f0bbbbbbb3)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefffffffffffff)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cf0ffcf0ffff)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffcffffffffff)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030fcfc3030)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdffffff)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff0008)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000030003)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500000005000000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00000f1f0000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf222f222f222f222)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff444f444)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c0000ffff00ff)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc4000ffff5000)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(LIOB33_X0Y155_IOB_X0Y155_I),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I2(1'b1),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000002)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcccccc5500f0f0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffefff55ff55ff)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfceefeeefe)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf555f0cc)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_A5Q),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0aaa0aee0eaa0a)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000ff2f2f2f2)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_AO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ff30ffbaffba)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cc00df53dc50)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba00babaaa00aaaa)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(LIOB33_X0Y153_IOB_X0Y153_I),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0fff0fff0f)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y153_IOB_X0Y153_I),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fafaaaaa)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I3(1'b1),
.I4(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f005f005f)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I1(1'b1),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b88b8b8888)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y122_SLICE_X18Y122_DO6),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff01fe00ff)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa3c00afaa0f00)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(LIOB33_X0Y161_IOB_X0Y161_I),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa5aaaa33363333)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1b1b100ff00ff)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.I2(CLBLM_R_X13Y122_SLICE_X19Y122_DO6),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0c0c)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.I1(CLBLM_R_X13Y122_SLICE_X19Y122_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8c83808fbcb3b0b)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_R_X13Y122_SLICE_X19Y122_DO6),
.I4(CLBLM_R_X15Y125_SLICE_X20Y125_BO6),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7e6b3a2d5c49180)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_DO6),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebadc9876325410)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0c0c0afa0cfcf)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e1f0e100010001)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h048c26ae159d37bf)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_BQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbea7362d9c85140)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_BQ),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaf0cc00aaf0cc)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.I1(CLBLM_R_X13Y122_SLICE_X19Y122_DO6),
.I2(CLBLM_R_X15Y125_SLICE_X20Y125_BO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0ffccaaf000cc)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I2(CLBLM_R_X15Y125_SLICE_X20Y125_BO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y122_SLICE_X19Y122_DO6),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0f33333333)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_CO6),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30eeeefc302222)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_CO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0eeee2222)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.I3(CLBLM_R_X13Y125_SLICE_X19Y125_CO6),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf3fa030af30a03)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_DO6),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_CO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeee4444)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_BO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_CO6),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h303f303f0505f5f5)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_R_X13Y127_SLICE_X19Y127_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000000000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff4fff444)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I1(LIOB33_X0Y155_IOB_X0Y155_I),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeffae55045504)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c44773f3f4477)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550f33ff550f33)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fcacaf000caca)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_R_X11Y125_SLICE_X14Y125_DO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfafc0a0cfa0c0a)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_DO6),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33aa33aa30a033aa)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffff00880000)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30ffffff)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(LIOB33_X0Y191_IOB_X0Y191_I),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I2(LIOB33_X0Y151_IOB_X0Y152_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330f0f33330f05)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550f0f55550f03)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_R_X15Y125_SLICE_X20Y125_DO6),
.I3(CLBLM_R_X15Y130_SLICE_X20Y130_BQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffff02000000)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefee33332322)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I3(LIOB33_X0Y155_IOB_X0Y156_I),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_AO6),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfefc3030ba30)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I5(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000010ffffff7f)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff40f0f0f04)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I1(LIOB33_X0Y155_IOB_X0Y155_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h500350035f035f03)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30053f0530f53ff5)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff10ff80)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeaf3c0f3c0f3c0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfafffffccaa)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.I5(LIOB33_X0Y157_IOB_X0Y157_I),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000004fffbffff)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ff8f80808)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_CO6),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f3535f0ff3535)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03f3505003f35f5f)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aeffae0c)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd0f0dfffc0f0c)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_BO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.I5(LIOB33_X0Y157_IOB_X0Y157_I),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h04c407c734f437f7)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffcfffafafcfc)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_DO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_DO6),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I5(LIOB33_X0Y155_IOB_X0Y155_I),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ff55e4e4aa00)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcacac0c0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I1(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_CO6),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd5fcc0fcc0fcc0f)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_CO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000000001)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ff22)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f3355000f3355ff)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500330f55ff330f)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a020a5f5f135f)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfcacfcfcfcfcf)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_BO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33550f0033550fff)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f3535f0ff3535)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50ffdcfffafffeff)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I1(LIOB33_X0Y151_IOB_X0Y151_I),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0cfc0cfcf)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_BO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fff000d0ddd00)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0fccee0faf)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf707f707ff0ff707)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_DO6),
.I1(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fff0ff404)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I1(LIOB33_X0Y151_IOB_X0Y152_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CO6),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X13Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f4fffff0f0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_DO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbfafaffbbfffa)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X13Y130_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I3(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fff30f03)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y130_SLICE_X13Y130_BO6),
.I4(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffffff)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffc30feba)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff808ff0ff808)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafa0a0acac)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(1'b1),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h03f303f30505f5f5)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I1(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h474747470033ccff)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff3fff0fff0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fffffff7f7)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff4f4ffffff44)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I1(LIOB33_X0Y155_IOB_X0Y155_I),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f0ff00)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I2(LIOB33_X0Y189_IOB_X0Y190_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfccffff0f003f33)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbb00110000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ffb0bfa0a)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X16Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X16Y100_DO5),
.O6(CLBLM_L_X12Y100_SLICE_X16Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X16Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X16Y100_CO5),
.O6(CLBLM_L_X12Y100_SLICE_X16Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X16Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X16Y100_BO5),
.O6(CLBLM_L_X12Y100_SLICE_X16Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X16Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X16Y100_AO5),
.O6(CLBLM_L_X12Y100_SLICE_X16Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X17Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X17Y100_DO5),
.O6(CLBLM_L_X12Y100_SLICE_X17Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X17Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X17Y100_CO5),
.O6(CLBLM_L_X12Y100_SLICE_X17Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y100_SLICE_X17Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y100_SLICE_X17Y100_BO5),
.O6(CLBLM_L_X12Y100_SLICE_X17Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000080000000)
  ) CLBLM_L_X12Y100_SLICE_X17Y100_ALUT (
.I0(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I1(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I4(CLBLM_R_X11Y102_SLICE_X14Y102_BO6),
.I5(CLBLM_L_X12Y102_SLICE_X17Y102_AO5),
.O5(CLBLM_L_X12Y100_SLICE_X17Y100_AO5),
.O6(CLBLM_L_X12Y100_SLICE_X17Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y101_SLICE_X16Y101_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y101_SLICE_X16Y101_BO6),
.Q(CLBLM_L_X12Y101_SLICE_X16Y101_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaafaaafaaafa)
  ) CLBLM_L_X12Y101_SLICE_X16Y101_DLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y101_SLICE_X14Y101_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_L_X12Y101_SLICE_X16Y101_DO5),
.O6(CLBLM_L_X12Y101_SLICE_X16Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0f0f08040a05)
  ) CLBLM_L_X12Y101_SLICE_X16Y101_CLUT (
.I0(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I2(CLBLM_L_X12Y103_SLICE_X16Y103_CO6),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_AO5),
.I4(CLBLM_R_X11Y101_SLICE_X15Y101_AO5),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_L_X12Y101_SLICE_X16Y101_CO5),
.O6(CLBLM_L_X12Y101_SLICE_X16Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcf8a8acfcfcfcf)
  ) CLBLM_L_X12Y101_SLICE_X16Y101_BLUT (
.I0(CLBLM_L_X12Y101_SLICE_X16Y101_DO6),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y102_SLICE_X15Y102_CO6),
.I5(CLBLM_L_X12Y101_SLICE_X16Y101_CO6),
.O5(CLBLM_L_X12Y101_SLICE_X16Y101_BO5),
.O6(CLBLM_L_X12Y101_SLICE_X16Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0080808080)
  ) CLBLM_L_X12Y101_SLICE_X16Y101_ALUT (
.I0(CLBLM_L_X10Y100_SLICE_X12Y100_BO6),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I3(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y101_SLICE_X16Y101_AO5),
.O6(CLBLM_L_X12Y101_SLICE_X16Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa003c3c3c3c)
  ) CLBLM_L_X12Y101_SLICE_X17Y101_DLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_BO6),
.I2(CLBLM_R_X11Y101_SLICE_X15Y101_AO6),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y101_SLICE_X17Y101_DO5),
.O6(CLBLM_L_X12Y101_SLICE_X17Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080800000000000)
  ) CLBLM_L_X12Y101_SLICE_X17Y101_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_CO6),
.I2(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_L_X12Y101_SLICE_X17Y101_DO6),
.I5(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.O5(CLBLM_L_X12Y101_SLICE_X17Y101_CO5),
.O6(CLBLM_L_X12Y101_SLICE_X17Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0880000000000000)
  ) CLBLM_L_X12Y101_SLICE_X17Y101_BLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I2(CLBLM_L_X12Y101_SLICE_X16Y101_AO6),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I5(CLBLM_R_X11Y101_SLICE_X14Y101_BO6),
.O5(CLBLM_L_X12Y101_SLICE_X17Y101_BO5),
.O6(CLBLM_L_X12Y101_SLICE_X17Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000080000000)
  ) CLBLM_L_X12Y101_SLICE_X17Y101_ALUT (
.I0(CLBLM_L_X10Y101_SLICE_X12Y101_BO6),
.I1(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I2(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I3(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.O5(CLBLM_L_X12Y101_SLICE_X17Y101_AO5),
.O6(CLBLM_L_X12Y101_SLICE_X17Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y102_SLICE_X16Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y102_SLICE_X16Y102_AO6),
.Q(CLBLM_L_X12Y102_SLICE_X16Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y102_SLICE_X16Y102_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y102_SLICE_X16Y102_BO6),
.Q(CLBLM_L_X12Y102_SLICE_X16Y102_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cc)
  ) CLBLM_L_X12Y102_SLICE_X16Y102_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y100_SLICE_X14Y100_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y102_SLICE_X16Y102_DO5),
.O6(CLBLM_L_X12Y102_SLICE_X16Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc5f550f00)
  ) CLBLM_L_X12Y102_SLICE_X16Y102_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_CO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_CO6),
.I4(CLBLM_R_X11Y102_SLICE_X15Y102_AO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y102_SLICE_X16Y102_CO5),
.O6(CLBLM_L_X12Y102_SLICE_X16Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffffffaa)
  ) CLBLM_L_X12Y102_SLICE_X16Y102_BLUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I3(CLBLM_R_X11Y101_SLICE_X15Y101_CO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_CO5),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y102_SLICE_X16Y102_BO5),
.O6(CLBLM_L_X12Y102_SLICE_X16Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0c0e0ffffccee)
  ) CLBLM_L_X12Y102_SLICE_X16Y102_ALUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_DO6),
.I1(CLBLM_R_X11Y102_SLICE_X14Y102_CO6),
.I2(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_R_X11Y103_SLICE_X15Y103_AO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y102_SLICE_X16Y102_AO5),
.O6(CLBLM_L_X12Y102_SLICE_X16Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4800000000000000)
  ) CLBLM_L_X12Y102_SLICE_X17Y102_DLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I2(CLBLM_R_X11Y102_SLICE_X14Y102_AO6),
.I3(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I4(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.O5(CLBLM_L_X12Y102_SLICE_X17Y102_DO5),
.O6(CLBLM_L_X12Y102_SLICE_X17Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h17e8ff00ff00ff00)
  ) CLBLM_L_X12Y102_SLICE_X17Y102_CLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I2(CLBLM_R_X11Y102_SLICE_X14Y102_AO6),
.I3(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I4(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.O5(CLBLM_L_X12Y102_SLICE_X17Y102_CO5),
.O6(CLBLM_L_X12Y102_SLICE_X17Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf078f078f0f0f0)
  ) CLBLM_L_X12Y102_SLICE_X17Y102_BLUT (
.I0(CLBLM_L_X10Y102_SLICE_X13Y102_CO6),
.I1(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I2(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.O5(CLBLM_L_X12Y102_SLICE_X17Y102_BO5),
.O6(CLBLM_L_X12Y102_SLICE_X17Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaaaa000000)
  ) CLBLM_L_X12Y102_SLICE_X17Y102_ALUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y102_SLICE_X17Y102_AO5),
.O6(CLBLM_L_X12Y102_SLICE_X17Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y103_SLICE_X16Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y103_SLICE_X16Y103_AO6),
.Q(CLBLM_L_X12Y103_SLICE_X16Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0f8f0f0e0f0e0)
  ) CLBLM_L_X12Y103_SLICE_X16Y103_DLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.O5(CLBLM_L_X12Y103_SLICE_X16Y103_DO5),
.O6(CLBLM_L_X12Y103_SLICE_X16Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f7080000ef10)
  ) CLBLM_L_X12Y103_SLICE_X16Y103_CLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.O5(CLBLM_L_X12Y103_SLICE_X16Y103_CO5),
.O6(CLBLM_L_X12Y103_SLICE_X16Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h090906060b040d02)
  ) CLBLM_L_X12Y103_SLICE_X16Y103_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y103_SLICE_X16Y103_BO5),
.O6(CLBLM_L_X12Y103_SLICE_X16Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff73ff730000ff73)
  ) CLBLM_L_X12Y103_SLICE_X16Y103_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I1(CLBLM_R_X11Y103_SLICE_X15Y103_CO6),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_DO6),
.I3(CLBLM_L_X12Y103_SLICE_X16Y103_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.O5(CLBLM_L_X12Y103_SLICE_X16Y103_AO5),
.O6(CLBLM_L_X12Y103_SLICE_X16Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y103_SLICE_X17Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y103_SLICE_X17Y103_AO6),
.Q(CLBLM_L_X12Y103_SLICE_X17Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c3003c00c3003c)
  ) CLBLM_L_X12Y103_SLICE_X17Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I2(CLBLM_L_X12Y103_SLICE_X16Y103_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y103_SLICE_X17Y103_DO5),
.O6(CLBLM_L_X12Y103_SLICE_X17Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000800000000000)
  ) CLBLM_L_X12Y103_SLICE_X17Y103_CLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I3(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I4(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I5(CLBLM_L_X10Y102_SLICE_X13Y102_CO6),
.O5(CLBLM_L_X12Y103_SLICE_X17Y103_CO5),
.O6(CLBLM_L_X12Y103_SLICE_X17Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaaaaaaaaaaaaa8)
  ) CLBLM_L_X12Y103_SLICE_X17Y103_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I5(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.O5(CLBLM_L_X12Y103_SLICE_X17Y103_BO5),
.O6(CLBLM_L_X12Y103_SLICE_X17Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffe00ee00fe)
  ) CLBLM_L_X12Y103_SLICE_X17Y103_ALUT (
.I0(CLBLM_L_X12Y103_SLICE_X17Y103_DO6),
.I1(CLBLM_R_X13Y103_SLICE_X18Y103_CO6),
.I2(CLBLM_L_X12Y102_SLICE_X17Y102_BO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.O5(CLBLM_L_X12Y103_SLICE_X17Y103_AO5),
.O6(CLBLM_L_X12Y103_SLICE_X17Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.Q(CLBLM_L_X12Y104_SLICE_X16Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.Q(CLBLM_L_X12Y104_SLICE_X16Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff8fffffff88)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_DLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I3(CLBLM_L_X12Y103_SLICE_X16Y103_BO5),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I5(CLBLM_L_X12Y101_SLICE_X17Y101_DO5),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_DO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff50dc)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I1(CLBLM_L_X12Y101_SLICE_X17Y101_DO5),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_DO6),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_CO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f0ccffe0f0eeff)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_BLUT (
.I0(CLBLM_R_X11Y101_SLICE_X14Y101_DO6),
.I1(CLBLM_L_X12Y103_SLICE_X16Y103_CO6),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I3(CLBLM_R_X11Y104_SLICE_X15Y104_AO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_BO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5b1f5f5f5a0)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I2(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I3(CLBLM_L_X12Y103_SLICE_X16Y103_BO5),
.I4(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_CO6),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_AO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_DO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_CO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_BO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_AO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b0a3b0ab3a0b3a0)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_CLUT (
.I0(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I1(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_BLUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I5(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbeeaaaafbfefafa)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_ALUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I2(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.I3(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0000005fa05fa0)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_ALUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I2(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I4(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000100)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cccc00cc00)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000000a)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f2f0f0f3)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_CLUT (
.I0(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeefeccfc)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_BLUT (
.I0(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I1(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff800078f078f0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I4(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000022222222)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I2(1'b1),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffb3ffffffa0)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_CLUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aa2800000a08)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I3(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaaafffffeee)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I3(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff44ffc7)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_DO6),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_AO5),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffebfffafffb)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.I1(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I2(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000f0ffff00ff)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_BO6),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0bbb0bbb0bbb0bb)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_ALUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_DO6),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_DO6),
.I2(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444444444444444)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000000ff0000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffcffddffcc)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I5(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafaaefbb)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_ALUT (
.I0(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_L_X12Y113_SLICE_X17Y113_CO6),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc35541ffc35541)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff950000ff95ff95)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f50000f5f5f5f5)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff5055f0ff5055)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d0c57035d0c5703)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I1(CLBLM_L_X12Y111_SLICE_X17Y111_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0ffe1fff0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ddee0d0e)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffff88ccaaff)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_DO6),
.I1(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X12Y112_SLICE_X17Y112_CO6),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeddeedd0000eedd)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1122222222222222)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0f99093303)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f002d00330099)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_ALUT (
.I0(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y111_SLICE_X17Y111_AO6),
.Q(CLBLM_L_X12Y111_SLICE_X17Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y111_SLICE_X17Y111_BO6),
.Q(CLBLM_L_X12Y111_SLICE_X17Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001010000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heedddddddddddddd)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcf4500cfcfcfcf)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X13Y110_SLICE_X18Y110_BO6),
.I5(CLBLM_L_X12Y111_SLICE_X17Y111_CO6),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf45cfcfcf00cfcf)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_CO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000010)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333336)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I3(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fafcfef0055ccdd)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_BLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_DO6),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_A5Q),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b0ffbbf0a0ffaa)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_ALUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X12Y112_SLICE_X16Y112_CO6),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fff80008000)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5775577503300330)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200ff00fd)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_ALUT (
.I0(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_AO5),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_AO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00660066f0f6f0f6)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_DLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_AO5),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88f88fff88f8f8f8)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_CLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f00f0f)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa33bbccee)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I4(CLBLM_L_X12Y113_SLICE_X17Y113_AO6),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_ALUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_AO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0eca0eca0eca0ec)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_A5Q),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f8f88ff8fff8888)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_BLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00abbababa)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_ALUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff507c507c507c)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_BO5),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff53ff7053537070)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdf505fdcfc50f0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_A5Q),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_BO6),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_DO6),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y115_SLICE_X17Y115_BO6),
.Q(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y115_SLICE_X17Y115_AO6),
.Q(CLBLM_L_X12Y115_SLICE_X17Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50737350ff73ff50)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.I4(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050cc000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_DO6),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_CO6),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa78f8)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_A5Q),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_BO6),
.I2(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y116_SLICE_X16Y116_AO5),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y116_SLICE_X16Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X16Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h773f7f33550f5f00)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_A5Q),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I5(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_L_X12Y116_SLICE_X16Y116_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_A5Q),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X16Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X16Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_AO5),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_AO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y116_SLICE_X17Y116_BO6),
.Q(CLBLM_L_X12Y116_SLICE_X17Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_DLUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I5(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_DO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444ff4ff44fff4)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_CLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_BO6),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_CO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f0000000)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_BO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLM_L_X12Y116_SLICE_X17Y116_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_CO6),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y116_SLICE_X17Y116_AO5),
.O6(CLBLM_L_X12Y116_SLICE_X17Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y117_SLICE_X16Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444f4f477ccf7fc)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AO5),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444f4f477ccf7fc)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_DO6),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I2(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaac000c000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_ALUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_DO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y117_SLICE_X17Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X17Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y117_SLICE_X17Y117_BO6),
.Q(CLBLM_L_X12Y117_SLICE_X17Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222ff22ff22)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_DLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3b3b3ffa0ffa0a0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_CLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I4(CLBLM_L_X12Y116_SLICE_X17Y116_BO5),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000abaeaeae)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_DO6),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaabe55550050)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_DO6),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X16Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f5b3a0)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(LIOB33_X0Y155_IOB_X0Y156_I),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcf8acf00)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I1(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y120_SLICE_X16Y120_BO6),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I5(CLBLM_L_X12Y120_SLICE_X16Y120_CO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000005)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff28ffffff00ffff)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5515555515555555)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0045454500004500)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X17Y121_DO6),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaeaeaeffaeff)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(LIOB33_X0Y153_IOB_X0Y153_I),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I4(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeeefafffafa)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafaf8caf00)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_CO6),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y121_SLICE_X17Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X17Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeaafafafefa)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555575)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I2(LIOB33_X0Y151_IOB_X0Y152_I),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff444f000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X12Y121_SLICE_X17Y121_CO6),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afacafa0afac)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y121_SLICE_X17Y121_BO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y122_SLICE_X16Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X16Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f330f33550055ff)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_DLUT (
.I0(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I1(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I2(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I4(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fff440f04)
  ) CLBLM_L_X12Y122_SLICE_X16Y122_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_DO6),
.I4(CLBLM_L_X12Y121_SLICE_X17Y121_AQ),
.I5(CLBLM_L_X12Y122_SLICE_X16Y122_CO6),
.O5(CLBLM_L_X12Y122_SLICE_X16Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X16Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y122_SLICE_X17Y122_AO6),
.Q(CLBLM_L_X12Y122_SLICE_X17Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_DO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000050)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_CLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I1(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I2(LIOB33_X0Y151_IOB_X0Y151_I),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_CO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff50730033)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I5(CLBLM_L_X12Y122_SLICE_X17Y122_CO6),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_BO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff30ff30)
  ) CLBLM_L_X12Y122_SLICE_X17Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I3(CLBLM_L_X12Y122_SLICE_X17Y122_BO6),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y122_SLICE_X17Y122_AO5),
.O6(CLBLM_L_X12Y122_SLICE_X17Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y123_SLICE_X16Y123_BO6),
.Q(CLBLM_L_X12Y123_SLICE_X16Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcffccffdc50cc00)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I1(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000001000000)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffa0aff0ffe0e)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_BLUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_DO6),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X15Y121_SLICE_X21Y121_AQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_CO5),
.I5(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ffcfe0c0e)
  ) CLBLM_L_X12Y123_SLICE_X16Y123_ALUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I5(CLBLM_L_X12Y127_SLICE_X16Y127_CO6),
.O5(CLBLM_L_X12Y123_SLICE_X16Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X16Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y123_SLICE_X17Y123_AO6),
.Q(CLBLM_L_X12Y123_SLICE_X17Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff303030ff30ff)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.I2(LIOB33_X0Y151_IOB_X0Y151_I),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I4(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_DO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff10ff40ff)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_DO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_CO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a003b333b33)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_BO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fafbfafb)
  ) CLBLM_L_X12Y123_SLICE_X17Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I2(CLBLM_L_X12Y122_SLICE_X17Y122_DO6),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y123_SLICE_X17Y123_AO5),
.O6(CLBLM_L_X12Y123_SLICE_X17Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y124_SLICE_X16Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X16Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedc7654ba983210)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h08194c5d2a3b6e7f)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I4(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f7f3c0c0d5c0)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0ccccfffa)
  ) CLBLM_L_X12Y124_SLICE_X16Y124_ALUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.I2(CLBLM_L_X12Y123_SLICE_X16Y123_CO6),
.I3(CLBLM_L_X12Y124_SLICE_X16Y124_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.O5(CLBLM_L_X12Y124_SLICE_X16Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X16Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y124_SLICE_X17Y124_AO6),
.Q(CLBLM_L_X12Y124_SLICE_X17Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h024613578ace9bdf)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_DO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd75b931ec64a820)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I5(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_CO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fff00dd00)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_BO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafacafafafacaf)
  ) CLBLM_L_X12Y124_SLICE_X17Y124_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X16Y123_BQ),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_BO6),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.O5(CLBLM_L_X12Y124_SLICE_X17Y124_AO5),
.O6(CLBLM_L_X12Y124_SLICE_X17Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_AO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y125_SLICE_X16Y125_BO6),
.Q(CLBLM_L_X12Y125_SLICE_X16Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ffe2e2e2)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I1(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10303030153f3f3f)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I2(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffddffcc)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_BLUT (
.I0(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.I2(CLBLM_L_X12Y125_SLICE_X16Y125_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_DO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007373ff00ffff)
  ) CLBLM_L_X12Y125_SLICE_X16Y125_ALUT (
.I0(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X12Y125_SLICE_X16Y125_CO6),
.O5(CLBLM_L_X12Y125_SLICE_X16Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X16Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h101310131c1f1c1f)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I4(1'b1),
.I5(CLBLM_R_X15Y125_SLICE_X21Y125_AQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_DO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00ff0f0f0077)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I3(CLBLM_R_X15Y125_SLICE_X20Y125_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X15Y129_SLICE_X20Y129_AQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_CO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00450055ff45ff55)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_BLUT (
.I0(CLBLM_L_X12Y125_SLICE_X17Y125_DO6),
.I1(CLBLM_R_X15Y127_SLICE_X20Y127_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_BO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h11110a5fbbbb0a5f)
  ) CLBLM_L_X12Y125_SLICE_X17Y125_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X15Y127_SLICE_X20Y127_AQ),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_R_X15Y125_SLICE_X21Y125_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.O5(CLBLM_L_X12Y125_SLICE_X17Y125_AO5),
.O6(CLBLM_L_X12Y125_SLICE_X17Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555505af05af)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0007f0ff7077)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008000ffbfffff)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1f5a0f5f5f5f5f5)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(CLBLM_L_X16Y126_SLICE_X22Y126_BO6),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_CO6),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y126_SLICE_X17Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X17Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004050c0d)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_DLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_AO6),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_CLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c3f04150c3f0c3f)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2ff020fffff0f0f)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_ALUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_BO6),
.I4(CLBLM_R_X15Y124_SLICE_X20Y124_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55fcf5cc55cc55)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I3(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000080)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff00dcdc)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_BLUT (
.I0(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_BO6),
.I2(LIOB33_X0Y151_IOB_X0Y152_I),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_AO6),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcacfcfcfcaca)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_ALUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_DO6),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.I5(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.Q(CLBLM_L_X12Y127_SLICE_X17Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaaffff0c005d55)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_DLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000100000)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ff0f30003)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I4(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_BO6),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcacacfca)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_ALUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I4(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfd5dfd5df)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_DLUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I1(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff33eca0ffb3)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I1(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffccafccaa)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_ALUT (
.I0(CLBLM_L_X12Y128_SLICE_X16Y128_DO6),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I2(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(CLBLM_L_X12Y128_SLICE_X16Y128_CO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y128_SLICE_X17Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X17Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff0ff33fff3)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcccc0fff00ff)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I2(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffab5501)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_BO6),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I5(CLBLM_L_X12Y128_SLICE_X17Y128_CO6),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafffafafafa)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I1(1'b1),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_DO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7f77772f2f2222)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_CLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I3(1'b1),
.I4(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004400000002)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0bbaa)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_ALUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_BO5),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000af8c0000af8c)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_DLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I4(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff03ffffffab)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_CLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I3(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.I4(CLBLM_L_X12Y129_SLICE_X17Y129_BO5),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000008000)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000002000)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88ffcc0a080f0c)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffc0f3eafb)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff33ff00)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_BO6),
.I4(LIOB33_X0Y151_IOB_X0Y152_I),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y130_SLICE_X17Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X17Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ffffff50ff50)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_CO6),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I5(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccdcccdcccdc)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I4(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa2222aaff2233)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X17Y130_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000000000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafabbbbfffaffbb)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffce3302ffce3302)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_ALUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(LIOB33_X0Y141_IOB_X0Y142_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X12Y131_SLICE_X17Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X17Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff377f055)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I4(LIOB33_X0Y151_IOB_X0Y152_I),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aafffa00fa)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y101_SLICE_X22Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y101_SLICE_X22Y101_AO6),
.Q(CLBLM_L_X16Y101_SLICE_X22Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h22ff222222ff2222)
  ) CLBLM_L_X16Y101_SLICE_X22Y101_DLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_BO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_CO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y101_SLICE_X22Y101_DO5),
.O6(CLBLM_L_X16Y101_SLICE_X22Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h57575d5d03030c0c)
  ) CLBLM_L_X16Y101_SLICE_X22Y101_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I1(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I3(1'b1),
.I4(CLBLM_L_X16Y101_SLICE_X22Y101_BO5),
.I5(CLBLM_L_X16Y102_SLICE_X22Y102_BO6),
.O5(CLBLM_L_X16Y101_SLICE_X22Y101_CO5),
.O6(CLBLM_L_X16Y101_SLICE_X22Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_L_X16Y101_SLICE_X22Y101_BLUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I1(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_CO6),
.I4(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y101_SLICE_X22Y101_BO5),
.O6(CLBLM_L_X16Y101_SLICE_X22Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3e2f3e2)
  ) CLBLM_L_X16Y101_SLICE_X22Y101_ALUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I3(CLBLM_R_X15Y103_SLICE_X21Y103_BO6),
.I4(1'b1),
.I5(CLBLM_L_X16Y101_SLICE_X22Y101_CO6),
.O5(CLBLM_L_X16Y101_SLICE_X22Y101_AO5),
.O6(CLBLM_L_X16Y101_SLICE_X22Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y101_SLICE_X23Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y101_SLICE_X23Y101_DO5),
.O6(CLBLM_L_X16Y101_SLICE_X23Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y101_SLICE_X23Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y101_SLICE_X23Y101_CO5),
.O6(CLBLM_L_X16Y101_SLICE_X23Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y101_SLICE_X23Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y101_SLICE_X23Y101_BO5),
.O6(CLBLM_L_X16Y101_SLICE_X23Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y101_SLICE_X23Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y101_SLICE_X23Y101_AO5),
.O6(CLBLM_L_X16Y101_SLICE_X23Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y102_SLICE_X22Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y102_SLICE_X22Y102_AO6),
.Q(CLBLM_L_X16Y102_SLICE_X22Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f030a020f030501)
  ) CLBLM_L_X16Y102_SLICE_X22Y102_DLUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_BO6),
.I1(CLBLM_L_X16Y102_SLICE_X23Y102_AO6),
.I2(CLBLM_R_X15Y103_SLICE_X21Y103_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I5(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.O5(CLBLM_L_X16Y102_SLICE_X22Y102_DO5),
.O6(CLBLM_L_X16Y102_SLICE_X22Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff0080000000)
  ) CLBLM_L_X16Y102_SLICE_X22Y102_CLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I2(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I3(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I4(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y102_SLICE_X22Y102_CO5),
.O6(CLBLM_L_X16Y102_SLICE_X22Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f078f080008000)
  ) CLBLM_L_X16Y102_SLICE_X22Y102_BLUT (
.I0(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I1(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y102_SLICE_X22Y102_BO5),
.O6(CLBLM_L_X16Y102_SLICE_X22Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd0ddd0ddd0ddd0d)
  ) CLBLM_L_X16Y102_SLICE_X22Y102_ALUT (
.I0(CLBLM_L_X16Y102_SLICE_X22Y102_DO6),
.I1(CLBLM_L_X16Y103_SLICE_X22Y103_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y102_SLICE_X22Y102_AO5),
.O6(CLBLM_L_X16Y102_SLICE_X22Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y102_SLICE_X23Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y102_SLICE_X23Y102_DO5),
.O6(CLBLM_L_X16Y102_SLICE_X23Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y102_SLICE_X23Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y102_SLICE_X23Y102_CO5),
.O6(CLBLM_L_X16Y102_SLICE_X23Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y102_SLICE_X23Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y102_SLICE_X23Y102_BO5),
.O6(CLBLM_L_X16Y102_SLICE_X23Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLM_L_X16Y102_SLICE_X23Y102_ALUT (
.I0(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I1(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I5(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.O5(CLBLM_L_X16Y102_SLICE_X23Y102_AO5),
.O6(CLBLM_L_X16Y102_SLICE_X23Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c3c300003c3c)
  ) CLBLM_L_X16Y103_SLICE_X22Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I2(CLBLM_R_X15Y103_SLICE_X21Y103_CO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_L_X16Y103_SLICE_X22Y103_DO5),
.O6(CLBLM_L_X16Y103_SLICE_X22Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h666c6ccc666c6ccc)
  ) CLBLM_L_X16Y103_SLICE_X22Y103_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I2(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X21Y100_CO6),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_CO5),
.I5(1'b1),
.O5(CLBLM_L_X16Y103_SLICE_X22Y103_CO5),
.O6(CLBLM_L_X16Y103_SLICE_X22Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdcffdcffdc)
  ) CLBLM_L_X16Y103_SLICE_X22Y103_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I1(CLBLM_L_X16Y103_SLICE_X23Y103_BO6),
.I2(CLBLM_R_X15Y103_SLICE_X20Y103_AO5),
.I3(CLBLM_R_X15Y103_SLICE_X21Y103_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X16Y103_SLICE_X22Y103_BO5),
.O6(CLBLM_L_X16Y103_SLICE_X22Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h090906063bcd37ce)
  ) CLBLM_L_X16Y103_SLICE_X22Y103_ALUT (
.I0(CLBLM_R_X15Y103_SLICE_X21Y103_CO6),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_R_X15Y102_SLICE_X21Y102_BO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_L_X16Y103_SLICE_X22Y103_AO5),
.O6(CLBLM_L_X16Y103_SLICE_X22Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h003caabe003caabe)
  ) CLBLM_L_X16Y103_SLICE_X23Y103_DLUT (
.I0(CLBLM_L_X16Y103_SLICE_X23Y103_AO6),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I2(CLBLM_R_X15Y100_SLICE_X21Y100_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y103_SLICE_X23Y103_DO5),
.O6(CLBLM_L_X16Y103_SLICE_X23Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X16Y103_SLICE_X23Y103_CLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I2(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I3(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I4(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I5(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.O5(CLBLM_L_X16Y103_SLICE_X23Y103_CO5),
.O6(CLBLM_L_X16Y103_SLICE_X23Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff888fffff8f88)
  ) CLBLM_L_X16Y103_SLICE_X23Y103_BLUT (
.I0(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_L_X16Y102_SLICE_X23Y102_AO6),
.I4(CLBLM_R_X15Y108_SLICE_X21Y108_AO6),
.I5(CLBLM_R_X15Y100_SLICE_X21Y100_CO6),
.O5(CLBLM_L_X16Y103_SLICE_X23Y103_BO5),
.O6(CLBLM_L_X16Y103_SLICE_X23Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_L_X16Y103_SLICE_X23Y103_ALUT (
.I0(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I2(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I3(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I4(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I5(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.O5(CLBLM_L_X16Y103_SLICE_X23Y103_AO5),
.O6(CLBLM_L_X16Y103_SLICE_X23Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y104_SLICE_X22Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y104_SLICE_X22Y104_AO6),
.Q(CLBLM_L_X16Y104_SLICE_X22Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y104_SLICE_X22Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y104_SLICE_X22Y104_BO6),
.Q(CLBLM_L_X16Y104_SLICE_X22Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1ef01ef078f078f0)
  ) CLBLM_L_X16Y104_SLICE_X22Y104_DLUT (
.I0(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I1(CLBLM_L_X16Y102_SLICE_X22Y102_BO5),
.I2(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I3(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I4(1'b1),
.I5(CLBLM_R_X15Y103_SLICE_X20Y103_DO6),
.O5(CLBLM_L_X16Y104_SLICE_X22Y104_DO5),
.O6(CLBLM_L_X16Y104_SLICE_X22Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000e0ee0000b0bb)
  ) CLBLM_L_X16Y104_SLICE_X22Y104_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I1(CLBLM_R_X15Y100_SLICE_X21Y100_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I3(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I4(CLBLM_L_X16Y108_SLICE_X22Y108_DO6),
.I5(CLBLM_L_X16Y102_SLICE_X23Y102_AO6),
.O5(CLBLM_L_X16Y104_SLICE_X22Y104_CO5),
.O6(CLBLM_L_X16Y104_SLICE_X22Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff3055555510)
  ) CLBLM_L_X16Y104_SLICE_X22Y104_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_L_X16Y104_SLICE_X22Y104_DO6),
.I3(CLBLM_R_X15Y105_SLICE_X20Y105_DO6),
.I4(CLBLM_L_X16Y103_SLICE_X22Y103_AO6),
.I5(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.O5(CLBLM_L_X16Y104_SLICE_X22Y104_BO5),
.O6(CLBLM_L_X16Y104_SLICE_X22Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550c04ff55ff55)
  ) CLBLM_L_X16Y104_SLICE_X22Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_DO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I4(CLBLM_L_X16Y103_SLICE_X22Y103_DO6),
.I5(CLBLM_R_X15Y104_SLICE_X21Y104_DO6),
.O5(CLBLM_L_X16Y104_SLICE_X22Y104_AO5),
.O6(CLBLM_L_X16Y104_SLICE_X22Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y104_SLICE_X23Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y104_SLICE_X23Y104_AO6),
.Q(CLBLM_L_X16Y104_SLICE_X23Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800800000000000)
  ) CLBLM_L_X16Y104_SLICE_X23Y104_DLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_CO6),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I2(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I3(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_CO5),
.I5(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.O5(CLBLM_L_X16Y104_SLICE_X23Y104_DO5),
.O6(CLBLM_L_X16Y104_SLICE_X23Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c7878f0f0f0f0f0)
  ) CLBLM_L_X16Y104_SLICE_X23Y104_CLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_CO6),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I2(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I3(CLBLM_L_X16Y102_SLICE_X22Y102_CO5),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I5(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.O5(CLBLM_L_X16Y104_SLICE_X23Y104_CO5),
.O6(CLBLM_L_X16Y104_SLICE_X23Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habffababbaffbaba)
  ) CLBLM_L_X16Y104_SLICE_X23Y104_BLUT (
.I0(CLBLM_L_X16Y103_SLICE_X23Y103_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I2(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLM_L_X16Y105_SLICE_X23Y105_AO6),
.I5(CLBLM_L_X16Y103_SLICE_X23Y103_CO6),
.O5(CLBLM_L_X16Y104_SLICE_X23Y104_BO5),
.O6(CLBLM_L_X16Y104_SLICE_X23Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5a0f5a0)
  ) CLBLM_L_X16Y104_SLICE_X23Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(1'b1),
.I2(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I3(CLBLM_L_X16Y104_SLICE_X23Y104_BO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y106_SLICE_X20Y106_CO6),
.O5(CLBLM_L_X16Y104_SLICE_X23Y104_AO5),
.O6(CLBLM_L_X16Y104_SLICE_X23Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y105_SLICE_X22Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y105_SLICE_X22Y105_AO6),
.Q(CLBLM_L_X16Y105_SLICE_X22Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa0055005500aa)
  ) CLBLM_L_X16Y105_SLICE_X22Y105_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_R_X15Y105_SLICE_X20Y105_CO6),
.I5(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.O5(CLBLM_L_X16Y105_SLICE_X22Y105_DO5),
.O6(CLBLM_L_X16Y105_SLICE_X22Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff4ffffff44)
  ) CLBLM_L_X16Y105_SLICE_X22Y105_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_L_X16Y105_SLICE_X23Y105_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(CLBLM_L_X16Y110_SLICE_X22Y110_DO6),
.I4(CLBLM_L_X16Y105_SLICE_X22Y105_DO6),
.I5(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.O5(CLBLM_L_X16Y105_SLICE_X22Y105_CO5),
.O6(CLBLM_L_X16Y105_SLICE_X22Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffaafffbfffa)
  ) CLBLM_L_X16Y105_SLICE_X22Y105_BLUT (
.I0(CLBLM_L_X16Y108_SLICE_X22Y108_AO5),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I3(CLBLM_L_X16Y110_SLICE_X22Y110_DO6),
.I4(CLBLM_L_X16Y105_SLICE_X23Y105_CO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_L_X16Y105_SLICE_X22Y105_BO5),
.O6(CLBLM_L_X16Y105_SLICE_X22Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffaaffee)
  ) CLBLM_L_X16Y105_SLICE_X22Y105_ALUT (
.I0(CLBLM_L_X16Y105_SLICE_X22Y105_DO6),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_CO6),
.I2(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I3(CLBLM_L_X16Y105_SLICE_X22Y105_BO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X16Y105_SLICE_X22Y105_AO5),
.O6(CLBLM_L_X16Y105_SLICE_X22Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080800000000000)
  ) CLBLM_L_X16Y105_SLICE_X23Y105_DLUT (
.I0(CLBLM_R_X15Y103_SLICE_X20Y103_DO6),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I2(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I3(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_BO5),
.I5(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.O5(CLBLM_L_X16Y105_SLICE_X23Y105_DO5),
.O6(CLBLM_L_X16Y105_SLICE_X23Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc6ccc6ccccccc)
  ) CLBLM_L_X16Y105_SLICE_X23Y105_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I1(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I2(CLBLM_L_X16Y102_SLICE_X22Y102_BO5),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I5(CLBLM_R_X15Y103_SLICE_X20Y103_DO6),
.O5(CLBLM_L_X16Y105_SLICE_X23Y105_CO5),
.O6(CLBLM_L_X16Y105_SLICE_X23Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080800000000000)
  ) CLBLM_L_X16Y105_SLICE_X23Y105_BLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_DO6),
.I1(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I2(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I3(CLBLM_L_X16Y103_SLICE_X23Y103_CO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.O5(CLBLM_L_X16Y105_SLICE_X23Y105_BO5),
.O6(CLBLM_L_X16Y105_SLICE_X23Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5555aacc000000)
  ) CLBLM_L_X16Y105_SLICE_X23Y105_ALUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_DO6),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I2(1'b1),
.I3(CLBLM_L_X16Y103_SLICE_X23Y103_CO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y105_SLICE_X23Y105_AO5),
.O6(CLBLM_L_X16Y105_SLICE_X23Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y106_SLICE_X22Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y106_SLICE_X22Y106_AO6),
.Q(CLBLM_L_X16Y106_SLICE_X22Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_L_X16Y106_SLICE_X22Y106_DLUT (
.I0(CLBLM_R_X15Y102_SLICE_X21Y102_BO6),
.I1(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I2(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I4(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I5(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.O5(CLBLM_L_X16Y106_SLICE_X22Y106_DO5),
.O6(CLBLM_L_X16Y106_SLICE_X22Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h15ff151540ff4040)
  ) CLBLM_L_X16Y106_SLICE_X22Y106_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I2(CLBLM_L_X16Y106_SLICE_X23Y106_BO5),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(CLBLM_L_X16Y106_SLICE_X22Y106_DO6),
.I5(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.O5(CLBLM_L_X16Y106_SLICE_X22Y106_CO5),
.O6(CLBLM_L_X16Y106_SLICE_X22Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc0ff006aaaaaaa)
  ) CLBLM_L_X16Y106_SLICE_X22Y106_BLUT (
.I0(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I1(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I2(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I3(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I4(CLBLM_R_X15Y102_SLICE_X21Y102_BO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y106_SLICE_X22Y106_BO5),
.O6(CLBLM_L_X16Y106_SLICE_X22Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbbbbbb8b8)
  ) CLBLM_L_X16Y106_SLICE_X22Y106_ALUT (
.I0(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y106_SLICE_X23Y106_CO6),
.I3(1'b1),
.I4(CLBLM_L_X16Y106_SLICE_X22Y106_CO6),
.I5(CLBLM_R_X15Y106_SLICE_X21Y106_DO6),
.O5(CLBLM_L_X16Y106_SLICE_X22Y106_AO5),
.O6(CLBLM_L_X16Y106_SLICE_X22Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00ff00ff00)
  ) CLBLM_L_X16Y106_SLICE_X23Y106_DLUT (
.I0(CLBLM_L_X16Y103_SLICE_X23Y103_CO6),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I2(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I3(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.O5(CLBLM_L_X16Y106_SLICE_X23Y106_DO5),
.O6(CLBLM_L_X16Y106_SLICE_X23Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h132017fa13205fa0)
  ) CLBLM_L_X16Y106_SLICE_X23Y106_CLUT (
.I0(CLBLM_L_X16Y106_SLICE_X23Y106_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I2(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I3(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I5(CLBLM_L_X16Y105_SLICE_X23Y105_BO6),
.O5(CLBLM_L_X16Y106_SLICE_X23Y106_CO5),
.O6(CLBLM_L_X16Y106_SLICE_X23Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000080000000)
  ) CLBLM_L_X16Y106_SLICE_X23Y106_BLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_AO6),
.I1(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I2(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I4(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y106_SLICE_X23Y106_BO5),
.O6(CLBLM_L_X16Y106_SLICE_X23Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000006ccccccc)
  ) CLBLM_L_X16Y106_SLICE_X23Y106_ALUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I1(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I2(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I3(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I4(CLBLM_L_X16Y103_SLICE_X23Y103_CO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y106_SLICE_X23Y106_AO5),
.O6(CLBLM_L_X16Y106_SLICE_X23Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y107_SLICE_X22Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y107_SLICE_X22Y107_AO6),
.Q(CLBLM_L_X16Y107_SLICE_X22Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a55aa55a)
  ) CLBLM_L_X16Y107_SLICE_X22Y107_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(1'b1),
.I2(CLBLM_R_X15Y107_SLICE_X21Y107_AO5),
.I3(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLM_L_X16Y107_SLICE_X22Y107_DO5),
.O6(CLBLM_L_X16Y107_SLICE_X22Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabfbafababfbafa)
  ) CLBLM_L_X16Y107_SLICE_X22Y107_CLUT (
.I0(CLBLM_L_X16Y107_SLICE_X23Y107_BO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I2(CLBLM_L_X16Y106_SLICE_X23Y106_AO5),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_DO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y107_SLICE_X22Y107_CO5),
.O6(CLBLM_L_X16Y107_SLICE_X22Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cf8a0000cf45)
  ) CLBLM_L_X16Y107_SLICE_X22Y107_BLUT (
.I0(CLBLM_L_X16Y104_SLICE_X23Y104_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I4(CLBLM_L_X16Y108_SLICE_X23Y108_AO6),
.I5(CLBLM_L_X16Y106_SLICE_X23Y106_AO5),
.O5(CLBLM_L_X16Y107_SLICE_X22Y107_BO5),
.O6(CLBLM_L_X16Y107_SLICE_X22Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f0e0f0aaffeeff)
  ) CLBLM_L_X16Y107_SLICE_X22Y107_ALUT (
.I0(CLBLM_L_X16Y107_SLICE_X22Y107_DO6),
.I1(CLBLM_L_X16Y107_SLICE_X23Y107_DO5),
.I2(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I3(CLBLM_L_X16Y107_SLICE_X22Y107_BO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X16Y107_SLICE_X22Y107_AO5),
.O6(CLBLM_L_X16Y107_SLICE_X22Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a33cc33cc)
  ) CLBLM_L_X16Y107_SLICE_X23Y107_DLUT (
.I0(CLBLM_L_X16Y105_SLICE_X23Y105_BO6),
.I1(CLBLM_L_X16Y106_SLICE_X22Y106_BO6),
.I2(CLBLM_L_X16Y106_SLICE_X23Y106_DO6),
.I3(CLBLM_L_X16Y105_SLICE_X23Y105_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y107_SLICE_X23Y107_DO5),
.O6(CLBLM_L_X16Y107_SLICE_X23Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03ab03ab0cae0cae)
  ) CLBLM_L_X16Y107_SLICE_X23Y107_CLUT (
.I0(CLBLM_L_X16Y106_SLICE_X22Y106_BO5),
.I1(CLBLM_L_X16Y106_SLICE_X23Y106_BO5),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.O5(CLBLM_L_X16Y107_SLICE_X23Y107_CO5),
.O6(CLBLM_L_X16Y107_SLICE_X23Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcdcddcdcdcdc)
  ) CLBLM_L_X16Y107_SLICE_X23Y107_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_BO6),
.I2(CLBLM_L_X16Y106_SLICE_X23Y106_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I5(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.O5(CLBLM_L_X16Y107_SLICE_X23Y107_BO5),
.O6(CLBLM_L_X16Y107_SLICE_X23Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33bb00aa)
  ) CLBLM_L_X16Y107_SLICE_X23Y107_ALUT (
.I0(CLBLM_L_X16Y106_SLICE_X23Y106_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLM_L_X16Y107_SLICE_X23Y107_DO6),
.I5(CLBLM_L_X16Y107_SLICE_X23Y107_CO6),
.O5(CLBLM_L_X16Y107_SLICE_X23Y107_AO5),
.O6(CLBLM_L_X16Y107_SLICE_X23Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y108_SLICE_X22Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y108_SLICE_X22Y108_BO6),
.Q(CLBLM_L_X16Y108_SLICE_X22Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4fff4f4f8fff8f8)
  ) CLBLM_L_X16Y108_SLICE_X22Y108_DLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y108_SLICE_X21Y108_AO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_R_X15Y110_SLICE_X21Y110_AO5),
.I5(CLBLM_R_X15Y108_SLICE_X20Y108_AO6),
.O5(CLBLM_L_X16Y108_SLICE_X22Y108_DO5),
.O6(CLBLM_L_X16Y108_SLICE_X22Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h21ff12ff21211212)
  ) CLBLM_L_X16Y108_SLICE_X22Y108_CLUT (
.I0(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X15Y107_SLICE_X21Y107_AO5),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(CLBLM_L_X16Y106_SLICE_X22Y106_BO6),
.O5(CLBLM_L_X16Y108_SLICE_X22Y108_CO5),
.O6(CLBLM_L_X16Y108_SLICE_X22Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55f351f050)
  ) CLBLM_L_X16Y108_SLICE_X22Y108_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_L_X16Y107_SLICE_X22Y107_CO6),
.I3(LIOB33_SING_X0Y149_IOB_X0Y149_I),
.I4(CLBLM_L_X16Y107_SLICE_X23Y107_DO5),
.I5(CLBLM_L_X16Y108_SLICE_X22Y108_CO6),
.O5(CLBLM_L_X16Y108_SLICE_X22Y108_BO5),
.O6(CLBLM_L_X16Y108_SLICE_X22Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00002f228f88)
  ) CLBLM_L_X16Y108_SLICE_X22Y108_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X16Y109_SLICE_X22Y109_BO6),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I3(CLBLM_L_X16Y109_SLICE_X22Y109_AO5),
.I4(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y108_SLICE_X22Y108_AO5),
.O6(CLBLM_L_X16Y108_SLICE_X22Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y108_SLICE_X23Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y108_SLICE_X23Y108_DO5),
.O6(CLBLM_L_X16Y108_SLICE_X23Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y108_SLICE_X23Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y108_SLICE_X23Y108_CO5),
.O6(CLBLM_L_X16Y108_SLICE_X23Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y108_SLICE_X23Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y108_SLICE_X23Y108_BO5),
.O6(CLBLM_L_X16Y108_SLICE_X23Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdffdcffcddddcccc)
  ) CLBLM_L_X16Y108_SLICE_X23Y108_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_BO6),
.I2(CLBLM_L_X16Y108_SLICE_X22Y108_AO6),
.I3(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I4(CLBLM_L_X16Y109_SLICE_X23Y109_AO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X16Y108_SLICE_X23Y108_AO5),
.O6(CLBLM_L_X16Y108_SLICE_X23Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f0f0f0f0f0)
  ) CLBLM_L_X16Y109_SLICE_X22Y109_DLUT (
.I0(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I2(CLBLM_R_X15Y107_SLICE_X21Y107_CQ),
.I3(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.I4(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I5(CLBLM_L_X16Y110_SLICE_X22Y110_BO6),
.O5(CLBLM_L_X16Y109_SLICE_X22Y109_DO5),
.O6(CLBLM_L_X16Y109_SLICE_X22Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00ff00ff00)
  ) CLBLM_L_X16Y109_SLICE_X22Y109_CLUT (
.I0(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I1(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I2(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I3(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I4(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I5(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.O5(CLBLM_L_X16Y109_SLICE_X22Y109_CO5),
.O6(CLBLM_L_X16Y109_SLICE_X22Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X16Y109_SLICE_X22Y109_BLUT (
.I0(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I3(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I4(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I5(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.O5(CLBLM_L_X16Y109_SLICE_X22Y109_BO5),
.O6(CLBLM_L_X16Y109_SLICE_X22Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a000003cf03cf0)
  ) CLBLM_L_X16Y109_SLICE_X22Y109_ALUT (
.I0(CLBLM_L_X16Y109_SLICE_X22Y109_BO6),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I2(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I3(CLBLM_L_X16Y110_SLICE_X22Y110_BO6),
.I4(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y109_SLICE_X22Y109_AO5),
.O6(CLBLM_L_X16Y109_SLICE_X22Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y109_SLICE_X23Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y109_SLICE_X23Y109_DO5),
.O6(CLBLM_L_X16Y109_SLICE_X23Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_L_X16Y109_SLICE_X23Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I4(1'b1),
.I5(CLBLM_L_X16Y110_SLICE_X22Y110_BO6),
.O5(CLBLM_L_X16Y109_SLICE_X23Y109_CO5),
.O6(CLBLM_L_X16Y109_SLICE_X23Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f1f0f0f0f0)
  ) CLBLM_L_X16Y109_SLICE_X23Y109_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.O5(CLBLM_L_X16Y109_SLICE_X23Y109_BO5),
.O6(CLBLM_L_X16Y109_SLICE_X23Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7878f0f07f80ff00)
  ) CLBLM_L_X16Y109_SLICE_X23Y109_ALUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I1(CLBLM_L_X16Y110_SLICE_X22Y110_BO6),
.I2(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I3(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.I4(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y109_SLICE_X23Y109_AO5),
.O6(CLBLM_L_X16Y109_SLICE_X23Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y110_SLICE_X22Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y110_SLICE_X22Y110_AO6),
.Q(CLBLM_L_X16Y110_SLICE_X22Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000030)
  ) CLBLM_L_X16Y110_SLICE_X22Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_L_X16Y110_SLICE_X22Y110_DO5),
.O6(CLBLM_L_X16Y110_SLICE_X22Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff8f888f88)
  ) CLBLM_L_X16Y110_SLICE_X22Y110_CLUT (
.I0(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_L_X16Y109_SLICE_X22Y109_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X16Y110_SLICE_X22Y110_CO5),
.O6(CLBLM_L_X16Y110_SLICE_X22Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X16Y110_SLICE_X22Y110_BLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I3(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I4(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I5(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.O5(CLBLM_L_X16Y110_SLICE_X22Y110_BO5),
.O6(CLBLM_L_X16Y110_SLICE_X22Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff4ff0000f4ff)
  ) CLBLM_L_X16Y110_SLICE_X22Y110_ALUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I1(CLBLM_L_X16Y109_SLICE_X22Y109_CO6),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO6),
.I3(CLBLM_R_X15Y111_SLICE_X20Y111_DO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.O5(CLBLM_L_X16Y110_SLICE_X22Y110_AO5),
.O6(CLBLM_L_X16Y110_SLICE_X22Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001100)
  ) CLBLM_L_X16Y110_SLICE_X23Y110_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_L_X16Y110_SLICE_X23Y110_DO5),
.O6(CLBLM_L_X16Y110_SLICE_X23Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafffaaaaafafa)
  ) CLBLM_L_X16Y110_SLICE_X23Y110_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(1'b1),
.I2(CLBLM_L_X16Y109_SLICE_X23Y109_AO6),
.I3(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.O5(CLBLM_L_X16Y110_SLICE_X23Y110_CO5),
.O6(CLBLM_L_X16Y110_SLICE_X23Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccccccdc)
  ) CLBLM_L_X16Y110_SLICE_X23Y110_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_L_X16Y110_SLICE_X23Y110_BO5),
.O6(CLBLM_L_X16Y110_SLICE_X23Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000004400)
  ) CLBLM_L_X16Y110_SLICE_X23Y110_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.O6(CLBLM_L_X16Y110_SLICE_X23Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y111_SLICE_X22Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y111_SLICE_X22Y111_AO6),
.Q(CLBLM_L_X16Y111_SLICE_X22Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y111_SLICE_X22Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y111_SLICE_X22Y111_BO6),
.Q(CLBLM_L_X16Y111_SLICE_X22Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2222f22f)
  ) CLBLM_L_X16Y111_SLICE_X22Y111_DLUT (
.I0(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I2(CLBLM_L_X16Y111_SLICE_X23Y111_DO6),
.I3(CLBLM_L_X16Y109_SLICE_X22Y109_AO5),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_R_X15Y111_SLICE_X20Y111_AO6),
.O5(CLBLM_L_X16Y111_SLICE_X22Y111_DO5),
.O6(CLBLM_L_X16Y111_SLICE_X22Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00f099f9)
  ) CLBLM_L_X16Y111_SLICE_X22Y111_CLUT (
.I0(CLBLM_L_X16Y109_SLICE_X23Y109_AO6),
.I1(CLBLM_L_X16Y111_SLICE_X23Y111_CO6),
.I2(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_BO6),
.O5(CLBLM_L_X16Y111_SLICE_X22Y111_CO5),
.O6(CLBLM_L_X16Y111_SLICE_X22Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaffff32323333)
  ) CLBLM_L_X16Y111_SLICE_X22Y111_BLUT (
.I0(CLBLM_L_X16Y111_SLICE_X22Y111_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y110_SLICE_X22Y110_CO6),
.I3(1'b1),
.I4(CLBLM_R_X15Y112_SLICE_X20Y112_BO6),
.I5(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.O5(CLBLM_L_X16Y111_SLICE_X22Y111_BO5),
.O6(CLBLM_L_X16Y111_SLICE_X22Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf8acf8acf)
  ) CLBLM_L_X16Y111_SLICE_X22Y111_ALUT (
.I0(CLBLM_L_X16Y110_SLICE_X23Y110_CO6),
.I1(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X15Y112_SLICE_X20Y112_CO6),
.I4(1'b1),
.I5(CLBLM_L_X16Y111_SLICE_X22Y111_CO6),
.O5(CLBLM_L_X16Y111_SLICE_X22Y111_AO5),
.O6(CLBLM_L_X16Y111_SLICE_X22Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y111_SLICE_X23Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y111_SLICE_X23Y111_AO6),
.Q(CLBLM_L_X16Y111_SLICE_X23Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000480000004)
  ) CLBLM_L_X16Y111_SLICE_X23Y111_DLUT (
.I0(CLBLM_R_X15Y110_SLICE_X21Y110_BO5),
.I1(CLBLM_R_X15Y110_SLICE_X20Y110_AO5),
.I2(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I4(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y111_SLICE_X23Y111_DO5),
.O6(CLBLM_L_X16Y111_SLICE_X23Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000004)
  ) CLBLM_L_X16Y111_SLICE_X23Y111_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I1(CLBLM_R_X15Y110_SLICE_X20Y110_AO5),
.I2(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I3(CLBLM_R_X15Y110_SLICE_X21Y110_BO5),
.I4(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I5(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.O5(CLBLM_L_X16Y111_SLICE_X23Y111_CO5),
.O6(CLBLM_L_X16Y111_SLICE_X23Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000300)
  ) CLBLM_L_X16Y111_SLICE_X23Y111_BLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.O6(CLBLM_L_X16Y111_SLICE_X23Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff75ff75)
  ) CLBLM_L_X16Y111_SLICE_X23Y111_ALUT (
.I0(CLBLM_R_X15Y111_SLICE_X20Y111_BO6),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I2(CLBLM_R_X15Y110_SLICE_X21Y110_AO5),
.I3(CLBLM_L_X16Y111_SLICE_X23Y111_BO6),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X16Y111_SLICE_X23Y111_AO5),
.O6(CLBLM_L_X16Y111_SLICE_X23Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y113_SLICE_X22Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X22Y113_DO5),
.O6(CLBLM_L_X16Y113_SLICE_X22Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X16Y113_SLICE_X22Y113_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I2(CLBLM_R_X15Y114_SLICE_X21Y114_CO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X22Y113_CO5),
.O6(CLBLM_L_X16Y113_SLICE_X22Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c000fc00fc00)
  ) CLBLM_L_X16Y113_SLICE_X22Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X22Y113_BO5),
.O6(CLBLM_L_X16Y113_SLICE_X22Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80008000c800c800)
  ) CLBLM_L_X16Y113_SLICE_X22Y113_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X22Y113_AO5),
.O6(CLBLM_L_X16Y113_SLICE_X22Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y113_SLICE_X23Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X23Y113_DO5),
.O6(CLBLM_L_X16Y113_SLICE_X23Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y113_SLICE_X23Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X23Y113_CO5),
.O6(CLBLM_L_X16Y113_SLICE_X23Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y113_SLICE_X23Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X23Y113_BO5),
.O6(CLBLM_L_X16Y113_SLICE_X23Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y113_SLICE_X23Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y113_SLICE_X23Y113_AO5),
.O6(CLBLM_L_X16Y113_SLICE_X23Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y114_SLICE_X22Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y114_SLICE_X22Y114_AO6),
.Q(CLBLM_L_X16Y114_SLICE_X22Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc005acccc)
  ) CLBLM_L_X16Y114_SLICE_X22Y114_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I1(CLBLM_L_X16Y114_SLICE_X22Y114_AQ),
.I2(CLBLM_L_X16Y113_SLICE_X22Y113_AO5),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.O5(CLBLM_L_X16Y114_SLICE_X22Y114_DO5),
.O6(CLBLM_L_X16Y114_SLICE_X22Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0aaa3aaa3aaa0a)
  ) CLBLM_L_X16Y114_SLICE_X22Y114_CLUT (
.I0(CLBLM_L_X16Y114_SLICE_X23Y114_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I5(CLBLM_L_X16Y113_SLICE_X22Y113_CO6),
.O5(CLBLM_L_X16Y114_SLICE_X22Y114_CO5),
.O6(CLBLM_L_X16Y114_SLICE_X22Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c8000000)
  ) CLBLM_L_X16Y114_SLICE_X22Y114_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y114_SLICE_X22Y114_BO5),
.O6(CLBLM_L_X16Y114_SLICE_X22Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeefefee22232322)
  ) CLBLM_L_X16Y114_SLICE_X22Y114_ALUT (
.I0(CLBLM_L_X16Y114_SLICE_X22Y114_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I4(CLBLM_L_X16Y113_SLICE_X22Y113_BO6),
.I5(CLBLM_R_X15Y114_SLICE_X21Y114_AQ),
.O5(CLBLM_L_X16Y114_SLICE_X22Y114_AO5),
.O6(CLBLM_L_X16Y114_SLICE_X22Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y114_SLICE_X23Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y114_SLICE_X23Y114_AO6),
.Q(CLBLM_L_X16Y114_SLICE_X23Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y114_SLICE_X23Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y114_SLICE_X23Y114_BO6),
.Q(CLBLM_L_X16Y114_SLICE_X23Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b88b8aaaaaaaa)
  ) CLBLM_L_X16Y114_SLICE_X23Y114_DLUT (
.I0(CLBLM_L_X16Y114_SLICE_X23Y114_BQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_L_X16Y114_SLICE_X22Y114_BO5),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_L_X16Y114_SLICE_X23Y114_DO5),
.O6(CLBLM_L_X16Y114_SLICE_X23Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888baaaa88b8aaaa)
  ) CLBLM_L_X16Y114_SLICE_X23Y114_CLUT (
.I0(CLBLM_L_X16Y115_SLICE_X23Y115_BQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_L_X16Y113_SLICE_X22Y113_CO5),
.O5(CLBLM_L_X16Y114_SLICE_X23Y114_CO5),
.O6(CLBLM_L_X16Y114_SLICE_X23Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeffe22222332)
  ) CLBLM_L_X16Y114_SLICE_X23Y114_BLUT (
.I0(CLBLM_L_X16Y114_SLICE_X23Y114_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y113_SLICE_X22Y113_AO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_L_X16Y114_SLICE_X22Y114_AQ),
.O5(CLBLM_L_X16Y114_SLICE_X23Y114_BO5),
.O6(CLBLM_L_X16Y114_SLICE_X23Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fd31fc30fe32)
  ) CLBLM_L_X16Y114_SLICE_X23Y114_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y114_SLICE_X22Y114_CO6),
.I3(CLBLM_L_X16Y115_SLICE_X23Y115_BQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_R_X15Y114_SLICE_X21Y114_BO5),
.O5(CLBLM_L_X16Y114_SLICE_X23Y114_AO5),
.O6(CLBLM_L_X16Y114_SLICE_X23Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y115_SLICE_X22Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y115_SLICE_X22Y115_AO6),
.Q(CLBLM_L_X16Y115_SLICE_X22Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a000000000)
  ) CLBLM_L_X16Y115_SLICE_X22Y115_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y114_SLICE_X21Y114_CO6),
.O5(CLBLM_L_X16Y115_SLICE_X22Y115_DO5),
.O6(CLBLM_L_X16Y115_SLICE_X22Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a00deccf000fccc)
  ) CLBLM_L_X16Y115_SLICE_X22Y115_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_L_X16Y115_SLICE_X22Y115_AQ),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.I4(CLBLM_L_X16Y116_SLICE_X23Y116_DO6),
.I5(CLBLM_R_X15Y114_SLICE_X21Y114_CO6),
.O5(CLBLM_L_X16Y115_SLICE_X22Y115_CO5),
.O6(CLBLM_L_X16Y115_SLICE_X22Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X16Y115_SLICE_X22Y115_BLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I2(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I3(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.O5(CLBLM_L_X16Y115_SLICE_X22Y115_BO5),
.O6(CLBLM_L_X16Y115_SLICE_X22Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb888b88b8)
  ) CLBLM_L_X16Y115_SLICE_X22Y115_ALUT (
.I0(CLBLM_R_X15Y115_SLICE_X21Y115_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y115_SLICE_X21Y115_BO6),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I5(CLBLM_L_X16Y115_SLICE_X22Y115_CO6),
.O5(CLBLM_L_X16Y115_SLICE_X22Y115_AO5),
.O6(CLBLM_L_X16Y115_SLICE_X22Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y115_SLICE_X23Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y115_SLICE_X23Y115_AO6),
.Q(CLBLM_L_X16Y115_SLICE_X23Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y115_SLICE_X23Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y115_SLICE_X23Y115_BO6),
.Q(CLBLM_L_X16Y115_SLICE_X23Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888dd8cccccccc)
  ) CLBLM_L_X16Y115_SLICE_X23Y115_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_L_X16Y115_SLICE_X23Y115_AQ),
.I2(CLBLM_L_X16Y115_SLICE_X22Y115_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_L_X16Y115_SLICE_X23Y115_DO5),
.O6(CLBLM_L_X16Y115_SLICE_X23Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800aa00aa00)
  ) CLBLM_L_X16Y115_SLICE_X23Y115_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y115_SLICE_X21Y115_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y115_SLICE_X23Y115_CO5),
.O6(CLBLM_L_X16Y115_SLICE_X23Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0d1f3f3c0e2)
  ) CLBLM_L_X16Y115_SLICE_X23Y115_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y115_SLICE_X23Y115_AQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I4(CLBLM_L_X16Y114_SLICE_X23Y114_CO6),
.I5(CLBLM_L_X16Y115_SLICE_X23Y115_CO6),
.O5(CLBLM_L_X16Y115_SLICE_X23Y115_BO5),
.O6(CLBLM_L_X16Y115_SLICE_X23Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafbfbfa0a0b0b0a)
  ) CLBLM_L_X16Y115_SLICE_X23Y115_ALUT (
.I0(CLBLM_L_X16Y115_SLICE_X23Y115_DO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I4(CLBLM_L_X16Y115_SLICE_X23Y115_CO5),
.I5(CLBLM_L_X16Y115_SLICE_X22Y115_AQ),
.O5(CLBLM_L_X16Y115_SLICE_X23Y115_AO5),
.O6(CLBLM_L_X16Y115_SLICE_X23Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fcf0f0f66cc0000)
  ) CLBLM_L_X16Y116_SLICE_X22Y116_DLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I2(CLBLM_L_X16Y116_SLICE_X23Y116_DO6),
.I3(CLBLM_R_X15Y114_SLICE_X20Y114_DO6),
.I4(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.I5(CLBLM_L_X16Y116_SLICE_X23Y116_BQ),
.O5(CLBLM_L_X16Y116_SLICE_X22Y116_DO5),
.O6(CLBLM_L_X16Y116_SLICE_X22Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X16Y116_SLICE_X22Y116_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(CLBLM_R_X15Y113_SLICE_X21Y113_BO6),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y116_SLICE_X22Y116_CO5),
.O6(CLBLM_L_X16Y116_SLICE_X22Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000000c000c000)
  ) CLBLM_L_X16Y116_SLICE_X22Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y113_SLICE_X21Y113_BO6),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I4(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y116_SLICE_X22Y116_BO5),
.O6(CLBLM_L_X16Y116_SLICE_X22Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X16Y116_SLICE_X22Y116_ALUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I4(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y116_SLICE_X22Y116_AO5),
.O6(CLBLM_L_X16Y116_SLICE_X22Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y116_SLICE_X23Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y116_SLICE_X23Y116_AO6),
.Q(CLBLM_L_X16Y116_SLICE_X23Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y116_SLICE_X23Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y116_SLICE_X23Y116_BO6),
.Q(CLBLM_L_X16Y116_SLICE_X23Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505050505050)
  ) CLBLM_L_X16Y116_SLICE_X23Y116_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(1'b1),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y116_SLICE_X23Y116_DO5),
.O6(CLBLM_L_X16Y116_SLICE_X23Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbf0004bfbb0400)
  ) CLBLM_L_X16Y116_SLICE_X23Y116_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_R_X15Y114_SLICE_X20Y114_DO6),
.I4(CLBLM_L_X16Y116_SLICE_X23Y116_AQ),
.I5(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.O5(CLBLM_L_X16Y116_SLICE_X23Y116_CO5),
.O6(CLBLM_L_X16Y116_SLICE_X23Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffde33003312)
  ) CLBLM_L_X16Y116_SLICE_X23Y116_BLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I3(CLBLM_L_X16Y116_SLICE_X22Y116_DO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_L_X16Y116_SLICE_X23Y116_AQ),
.O5(CLBLM_L_X16Y116_SLICE_X23Y116_BO5),
.O6(CLBLM_L_X16Y116_SLICE_X23Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3c0c0d1e2)
  ) CLBLM_L_X16Y116_SLICE_X23Y116_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y114_SLICE_X23Y114_BQ),
.I3(CLBLM_L_X16Y114_SLICE_X22Y114_BO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_L_X16Y116_SLICE_X23Y116_CO6),
.O5(CLBLM_L_X16Y116_SLICE_X23Y116_AO5),
.O6(CLBLM_L_X16Y116_SLICE_X23Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y117_SLICE_X22Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y117_SLICE_X22Y117_AO6),
.Q(CLBLM_L_X16Y117_SLICE_X22Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y117_SLICE_X22Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y117_SLICE_X22Y117_BO6),
.Q(CLBLM_L_X16Y117_SLICE_X22Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0e4f0f0f0f0)
  ) CLBLM_L_X16Y117_SLICE_X22Y117_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_L_X16Y116_SLICE_X22Y116_CO6),
.I2(CLBLM_L_X16Y117_SLICE_X22Y117_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_L_X16Y117_SLICE_X22Y117_DO5),
.O6(CLBLM_L_X16Y117_SLICE_X22Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0e2f0f0f0f0)
  ) CLBLM_L_X16Y117_SLICE_X22Y117_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_L_X16Y117_SLICE_X22Y117_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_L_X16Y116_SLICE_X22Y116_CO5),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_L_X16Y117_SLICE_X22Y117_CO5),
.O6(CLBLM_L_X16Y117_SLICE_X22Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0bbf0bbf0aa)
  ) CLBLM_L_X16Y117_SLICE_X22Y117_BLUT (
.I0(CLBLM_L_X16Y117_SLICE_X22Y117_DO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I2(CLBLM_L_X16Y117_SLICE_X22Y117_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I5(CLBLM_L_X16Y116_SLICE_X22Y116_AO5),
.O5(CLBLM_L_X16Y117_SLICE_X22Y117_BO5),
.O6(CLBLM_L_X16Y117_SLICE_X22Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd888d8d88)
  ) CLBLM_L_X16Y117_SLICE_X22Y117_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X15Y116_SLICE_X21Y116_BQ),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I3(CLBLM_L_X16Y116_SLICE_X22Y116_BO6),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I5(CLBLM_L_X16Y117_SLICE_X22Y117_CO6),
.O5(CLBLM_L_X16Y117_SLICE_X22Y117_AO5),
.O6(CLBLM_L_X16Y117_SLICE_X22Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y117_SLICE_X23Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y117_SLICE_X23Y117_DO5),
.O6(CLBLM_L_X16Y117_SLICE_X23Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y117_SLICE_X23Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y117_SLICE_X23Y117_CO5),
.O6(CLBLM_L_X16Y117_SLICE_X23Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101ff00f202ff00)
  ) CLBLM_L_X16Y117_SLICE_X23Y117_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_L_X16Y117_SLICE_X23Y117_AO5),
.O5(CLBLM_L_X16Y117_SLICE_X23Y117_BO5),
.O6(CLBLM_L_X16Y117_SLICE_X23Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880088880000)
  ) CLBLM_L_X16Y117_SLICE_X23Y117_ALUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I2(1'b1),
.I3(CLBLM_L_X16Y115_SLICE_X22Y115_BO6),
.I4(CLBLM_R_X15Y115_SLICE_X21Y115_DO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y117_SLICE_X23Y117_AO5),
.O6(CLBLM_L_X16Y117_SLICE_X23Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y118_SLICE_X22Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y118_SLICE_X22Y118_DO5),
.O6(CLBLM_L_X16Y118_SLICE_X22Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y118_SLICE_X22Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y118_SLICE_X22Y118_CO5),
.O6(CLBLM_L_X16Y118_SLICE_X22Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y118_SLICE_X22Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y118_SLICE_X22Y118_BO5),
.O6(CLBLM_L_X16Y118_SLICE_X22Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X16Y118_SLICE_X22Y118_ALUT (
.I0(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I1(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I2(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I3(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I4(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I5(CLBLM_R_X15Y118_SLICE_X20Y118_DO6),
.O5(CLBLM_L_X16Y118_SLICE_X22Y118_AO5),
.O6(CLBLM_L_X16Y118_SLICE_X22Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y118_SLICE_X23Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y118_SLICE_X23Y118_AO6),
.Q(CLBLM_L_X16Y118_SLICE_X23Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y118_SLICE_X23Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y118_SLICE_X23Y118_DO5),
.O6(CLBLM_L_X16Y118_SLICE_X23Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a0a0a0a0)
  ) CLBLM_L_X16Y118_SLICE_X23Y118_CLUT (
.I0(CLBLM_R_X15Y115_SLICE_X21Y115_DO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y118_SLICE_X23Y118_CO5),
.O6(CLBLM_L_X16Y118_SLICE_X23Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1f0f0d1c0f0f0)
  ) CLBLM_L_X16Y118_SLICE_X23Y118_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_L_X16Y118_SLICE_X23Y118_AQ),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_L_X16Y118_SLICE_X23Y118_CO6),
.O5(CLBLM_L_X16Y118_SLICE_X23Y118_BO5),
.O6(CLBLM_L_X16Y118_SLICE_X23Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff5a)
  ) CLBLM_L_X16Y118_SLICE_X23Y118_ALUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I1(CLBLM_R_X15Y117_SLICE_X21Y117_BQ),
.I2(CLBLM_L_X16Y115_SLICE_X22Y115_BO6),
.I3(CLBLM_L_X16Y118_SLICE_X23Y118_BO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X16Y118_SLICE_X23Y118_AO5),
.O6(CLBLM_L_X16Y118_SLICE_X23Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y119_SLICE_X22Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y119_SLICE_X22Y119_AO6),
.Q(CLBLM_L_X16Y119_SLICE_X22Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0ccc0ccc5cccac)
  ) CLBLM_L_X16Y119_SLICE_X22Y119_DLUT (
.I0(CLBLM_L_X16Y119_SLICE_X22Y119_CO5),
.I1(CLBLM_L_X16Y119_SLICE_X22Y119_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_L_X16Y119_SLICE_X22Y119_DO5),
.O6(CLBLM_L_X16Y119_SLICE_X22Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_L_X16Y119_SLICE_X22Y119_CLUT (
.I0(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I1(CLBLM_R_X15Y118_SLICE_X20Y118_DO6),
.I2(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I3(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I4(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y119_SLICE_X22Y119_CO5),
.O6(CLBLM_L_X16Y119_SLICE_X22Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80808080c0c0c0c0)
  ) CLBLM_L_X16Y119_SLICE_X22Y119_BLUT (
.I0(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I1(CLBLM_R_X15Y117_SLICE_X21Y117_CO6),
.I2(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y119_SLICE_X22Y119_BO5),
.O6(CLBLM_L_X16Y119_SLICE_X22Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000abbaabba)
  ) CLBLM_L_X16Y119_SLICE_X22Y119_ALUT (
.I0(CLBLM_L_X16Y119_SLICE_X22Y119_DO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I3(CLBLM_L_X16Y119_SLICE_X22Y119_BO6),
.I4(CLBLM_L_X16Y119_SLICE_X23Y119_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_L_X16Y119_SLICE_X22Y119_AO5),
.O6(CLBLM_L_X16Y119_SLICE_X22Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y119_SLICE_X23Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y119_SLICE_X23Y119_AO6),
.Q(CLBLM_L_X16Y119_SLICE_X23Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y119_SLICE_X23Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y119_SLICE_X23Y119_DO5),
.O6(CLBLM_L_X16Y119_SLICE_X23Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y119_SLICE_X23Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y119_SLICE_X23Y119_CO5),
.O6(CLBLM_L_X16Y119_SLICE_X23Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf050f072f072f050)
  ) CLBLM_L_X16Y119_SLICE_X23Y119_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_L_X16Y119_SLICE_X23Y119_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I5(CLBLM_R_X15Y119_SLICE_X20Y119_BO6),
.O5(CLBLM_L_X16Y119_SLICE_X23Y119_BO5),
.O6(CLBLM_L_X16Y119_SLICE_X23Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcdffce33013302)
  ) CLBLM_L_X16Y119_SLICE_X23Y119_ALUT (
.I0(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I3(CLBLM_L_X16Y119_SLICE_X23Y119_BO6),
.I4(CLBLM_L_X16Y119_SLICE_X22Y119_BO5),
.I5(CLBLM_R_X15Y119_SLICE_X20Y119_AQ),
.O5(CLBLM_L_X16Y119_SLICE_X23Y119_AO5),
.O6(CLBLM_L_X16Y119_SLICE_X23Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y121_SLICE_X22Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y121_SLICE_X22Y121_AO6),
.Q(CLBLM_L_X16Y121_SLICE_X22Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X22Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X22Y121_DO5),
.O6(CLBLM_L_X16Y121_SLICE_X22Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X22Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X22Y121_CO5),
.O6(CLBLM_L_X16Y121_SLICE_X22Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X22Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X22Y121_BO5),
.O6(CLBLM_L_X16Y121_SLICE_X22Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaccaaffaafc)
  ) CLBLM_L_X16Y121_SLICE_X22Y121_ALUT (
.I0(CLBLM_R_X15Y122_SLICE_X20Y122_AQ),
.I1(CLBLM_L_X16Y123_SLICE_X22Y123_AO6),
.I2(LIOB33_X0Y155_IOB_X0Y155_I),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y121_SLICE_X21Y121_BO6),
.I5(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.O5(CLBLM_L_X16Y121_SLICE_X22Y121_AO5),
.O6(CLBLM_L_X16Y121_SLICE_X22Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X23Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X23Y121_DO5),
.O6(CLBLM_L_X16Y121_SLICE_X23Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X23Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X23Y121_CO5),
.O6(CLBLM_L_X16Y121_SLICE_X23Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X23Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X23Y121_BO5),
.O6(CLBLM_L_X16Y121_SLICE_X23Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y121_SLICE_X23Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y121_SLICE_X23Y121_AO5),
.O6(CLBLM_L_X16Y121_SLICE_X23Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y123_SLICE_X22Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X22Y123_DO5),
.O6(CLBLM_L_X16Y123_SLICE_X22Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y123_SLICE_X22Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X22Y123_CO5),
.O6(CLBLM_L_X16Y123_SLICE_X22Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccccccce)
  ) CLBLM_L_X16Y123_SLICE_X22Y123_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X15Y124_SLICE_X21Y124_DO6),
.O5(CLBLM_L_X16Y123_SLICE_X22Y123_BO5),
.O6(CLBLM_L_X16Y123_SLICE_X22Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00040000ff7fffff)
  ) CLBLM_L_X16Y123_SLICE_X22Y123_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X22Y123_AO5),
.O6(CLBLM_L_X16Y123_SLICE_X22Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y123_SLICE_X23Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X23Y123_DO5),
.O6(CLBLM_L_X16Y123_SLICE_X23Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y123_SLICE_X23Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X23Y123_CO5),
.O6(CLBLM_L_X16Y123_SLICE_X23Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y123_SLICE_X23Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X23Y123_BO5),
.O6(CLBLM_L_X16Y123_SLICE_X23Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y123_SLICE_X23Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y123_SLICE_X23Y123_AO5),
.O6(CLBLM_L_X16Y123_SLICE_X23Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y125_SLICE_X22Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y125_SLICE_X22Y125_AO6),
.Q(CLBLM_L_X16Y125_SLICE_X22Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcfefcfcfcfcf)
  ) CLBLM_L_X16Y125_SLICE_X22Y125_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I2(CLBLM_L_X16Y125_SLICE_X23Y125_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X16Y125_SLICE_X22Y125_DO5),
.O6(CLBLM_L_X16Y125_SLICE_X22Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfccafaaccccaaaa)
  ) CLBLM_L_X16Y125_SLICE_X22Y125_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_L_X16Y125_SLICE_X22Y125_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_L_X16Y125_SLICE_X22Y125_CO5),
.O6(CLBLM_L_X16Y125_SLICE_X22Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000dfffffff)
  ) CLBLM_L_X16Y125_SLICE_X22Y125_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y125_SLICE_X22Y125_BO5),
.O6(CLBLM_L_X16Y125_SLICE_X22Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafa0afafafac)
  ) CLBLM_L_X16Y125_SLICE_X22Y125_ALUT (
.I0(CLBLM_L_X16Y126_SLICE_X22Y126_AQ),
.I1(LIOB33_X0Y155_IOB_X0Y155_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X16Y125_SLICE_X22Y125_BO6),
.I4(CLBLM_L_X16Y125_SLICE_X22Y125_CO6),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.O5(CLBLM_L_X16Y125_SLICE_X22Y125_AO5),
.O6(CLBLM_L_X16Y125_SLICE_X22Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaabfbb0f003f33)
  ) CLBLM_L_X16Y125_SLICE_X23Y125_DLUT (
.I0(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X16Y125_SLICE_X23Y125_DO5),
.O6(CLBLM_L_X16Y125_SLICE_X23Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000b0000000b000b)
  ) CLBLM_L_X16Y125_SLICE_X23Y125_CLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I2(CLBLM_L_X16Y125_SLICE_X23Y125_AO5),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_AO6),
.O5(CLBLM_L_X16Y125_SLICE_X23Y125_CO5),
.O6(CLBLM_L_X16Y125_SLICE_X23Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555000001110)
  ) CLBLM_L_X16Y125_SLICE_X23Y125_BLUT (
.I0(CLBLM_R_X15Y127_SLICE_X21Y127_AO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I4(CLBLM_L_X16Y125_SLICE_X23Y125_AO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O5(CLBLM_L_X16Y125_SLICE_X23Y125_BO5),
.O6(CLBLM_L_X16Y125_SLICE_X23Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000002000)
  ) CLBLM_L_X16Y125_SLICE_X23Y125_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y125_SLICE_X23Y125_AO5),
.O6(CLBLM_L_X16Y125_SLICE_X23Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y126_SLICE_X22Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_L_X16Y126_SLICE_X22Y126_AO6),
.Q(CLBLM_L_X16Y126_SLICE_X22Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLM_L_X16Y126_SLICE_X22Y126_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.O5(CLBLM_L_X16Y126_SLICE_X22Y126_DO5),
.O6(CLBLM_L_X16Y126_SLICE_X22Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfefffffc0ea)
  ) CLBLM_L_X16Y126_SLICE_X22Y126_CLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_L_X16Y126_SLICE_X22Y126_AQ),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.I4(CLBLM_L_X16Y126_SLICE_X22Y126_DO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_L_X16Y126_SLICE_X22Y126_CO5),
.O6(CLBLM_L_X16Y126_SLICE_X22Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffff00004000)
  ) CLBLM_L_X16Y126_SLICE_X22Y126_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y126_SLICE_X22Y126_BO5),
.O6(CLBLM_L_X16Y126_SLICE_X22Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff003030)
  ) CLBLM_L_X16Y126_SLICE_X22Y126_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(CLBLM_R_X13Y124_SLICE_X18Y124_BQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X16Y126_SLICE_X22Y126_CO6),
.O5(CLBLM_L_X16Y126_SLICE_X22Y126_AO5),
.O6(CLBLM_L_X16Y126_SLICE_X22Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y126_SLICE_X23Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y126_SLICE_X23Y126_DO5),
.O6(CLBLM_L_X16Y126_SLICE_X23Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033110301)
  ) CLBLM_L_X16Y126_SLICE_X23Y126_CLUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_AO6),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_BO6),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_AO5),
.O5(CLBLM_L_X16Y126_SLICE_X23Y126_CO5),
.O6(CLBLM_L_X16Y126_SLICE_X23Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5ffff5fffffff)
  ) CLBLM_L_X16Y126_SLICE_X23Y126_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.O6(CLBLM_L_X16Y126_SLICE_X23Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000a00000000a)
  ) CLBLM_L_X16Y126_SLICE_X23Y126_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.O6(CLBLM_L_X16Y126_SLICE_X23Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb22bb22bb2222)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf0f0f0aa0055ff)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h336633cc88000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaafc30fc30)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_A5Q),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcff303fcccf000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd8d8df8f88888)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_A5Q),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_A5Q),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaccffeeaacc00)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccff0ffcccf000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefc5c5eaeac0c0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f5a0f5a0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h555555551d1d1d1d)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550000ff55ff55)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff4ffff4444)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff00ccccffff)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcfefcfeecceecc)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0031313100313131)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30001000ffff5555)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(LIOB33_X0Y161_IOB_X0Y162_I),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb0baa0aaa0aaa0a)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(LIOB33_X0Y153_IOB_X0Y154_I),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdc50ffffdc50)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h007f00ff00ff00ff)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff5530100000)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(LIOB33_X0Y151_IOB_X0Y151_I),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffc8888888)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000580000000)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffea00aa00ea)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I1(LIOB33_X0Y161_IOB_X0Y161_I),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I5(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X2Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00aaaaffaa)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(LIOB33_X0Y151_IOB_X0Y151_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0aff0aff0a)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555dff7f00cc00cc)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f022ff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeeafaaefeeafaa)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafe00cc0ace00cc)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(LIOB33_X0Y151_IOB_X0Y152_I),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0aaaae0a0eeaa)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(LIOB33_X0Y155_IOB_X0Y155_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafaf23af00)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I4(LIOB33_X0Y151_IOB_X0Y152_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdcffdcdcdcdcdc)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacac0000ffacff00)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I1(LIOB33_X0Y153_IOB_X0Y153_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaea0000aaeaaaea)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I1(LIOB33_X0Y155_IOB_X0Y156_I),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a8a8acfcfcfcf)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ff444444ff4444)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(LIOB33_X0Y159_IOB_X0Y160_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcceecceecceecc)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffccff00ff00)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000077773f77)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(LIOB33_X0Y159_IOB_X0Y160_I),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I3(LIOB33_X0Y185_IOB_X0Y185_I),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h37df135d5d454504)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcffffffff)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5d4e8a0d450f5d4)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5ddf5d45044504)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000696600009699)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he800fe80ffe8b332)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00f0000cccc)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h07fff800ffff0000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000007fff8000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc55aaddee)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.I2(1'b1),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f9f0f6f00990066)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeaa880fcc0fcc0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000036cc66cc)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5d4504cf0ccf0c)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I4(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00f53707053)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ffe0efe0e)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050a0a0a0a0505)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2211221111221122)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbffe3bbc23380220)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000100010001fffe)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6339399c9cc6c663)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafefafffffefa)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc936996636c96699)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fca800a00f000f0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4114ffffc33c)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h030c030c339dcf6e)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000004b2db4d2)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fffffa00fa)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa5555aa55aa)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550faf00550faf)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0013cc7f11017737)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h996639c6cc339c63)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccfcc0f000f00)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f00030f0f0303)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaf0eef0aa)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(LIOB33_X0Y163_IOB_X0Y164_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00800088f0f0ffff)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(LIOB33_X0Y157_IOB_X0Y158_I),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff03f3ffff)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y157_IOB_X0Y158_I),
.I2(LIOB33_X0Y185_IOB_X0Y185_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000b080ff00ff80)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(LIOB33_X0Y163_IOB_X0Y164_I),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fa32fa32fa32)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fdfdfdfd)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h330033003300ff00)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I4(LIOB33_X0Y185_IOB_X0Y185_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f300f033f300f0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0133013303330333)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ff3133f0ff3033)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a000a000a000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y159_IOB_X0Y159_I),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0f0f000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb0ab300bb00bb00)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(LIOB33_X0Y163_IOB_X0Y163_I),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0307030707070707)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc8000cccc0000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaf0aafc)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffefe)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000008880000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.I2(LIOB33_X0Y185_IOB_X0Y185_I),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefeee0000feee)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffb000000000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004fffbffff0000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeaaaaaaaaaaa)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50ae04fe54)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X13Y118_SLICE_X18Y118_AO6),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I4(LIOB33_X0Y181_IOB_X0Y182_I),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_BO6),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa0f0afffc0f0c)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(LIOB33_X0Y181_IOB_X0Y182_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BO6),
.I4(LIOB33_X0Y197_IOB_X0Y198_I),
.I5(CLBLM_R_X13Y118_SLICE_X18Y118_AO6),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0a0bbaae0a0eeaa)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff007f7f8080)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffccccfa50)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(CLBLM_R_X13Y118_SLICE_X18Y118_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(LIOB33_X0Y181_IOB_X0Y182_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_BO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500550055)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddccccffccffcc)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I4(LIOB33_X0Y163_IOB_X0Y163_I),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c0c0c0c0c0c0c0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffc0f0d0f0c)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.I4(LIOB33_X0Y177_IOB_X0Y178_I),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f0f033330000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I5(LIOB33_X0Y161_IOB_X0Y162_I),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011005555555555)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaa0e0affff0f0f)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fa00aaf0fa00aa)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(LIOB33_X0Y179_IOB_X0Y180_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafaaafaaafaaa)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fbbaa0b0a)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_X0Y177_IOB_X0Y177_I),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc50dc50dc50dc50)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(LIOB33_X0Y179_IOB_X0Y179_I),
.I3(LIOB33_X0Y163_IOB_X0Y163_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fcf0fcf0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I3(LIOB33_X0Y159_IOB_X0Y160_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaf0ffff0000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0faaee0a0e)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.I1(LIOB33_X0Y175_IOB_X0Y176_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(LIOB33_X0Y163_IOB_X0Y163_I),
.I1(1'b1),
.I2(LIOB33_X0Y165_IOB_X0Y165_I),
.I3(1'b1),
.I4(LIOB33_X0Y163_IOB_X0Y164_I),
.I5(LIOB33_X0Y151_IOB_X0Y151_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y153_I),
.I1(LIOB33_X0Y155_IOB_X0Y155_I),
.I2(LIOB33_X0Y151_IOB_X0Y152_I),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.I4(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.I5(LIOB33_X0Y153_IOB_X0Y154_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003c2c3c3c)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(LIOB33_X0Y183_IOB_X0Y183_I),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(LIOB33_X0Y183_IOB_X0Y184_I),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff3f0000ff7f)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(LIOB33_X0Y183_IOB_X0Y183_I),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf0ffffd8100000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I2(LIOB33_X0Y183_IOB_X0Y183_I),
.I3(LIOB33_X0Y185_IOB_X0Y185_I),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccbf00cf00)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I2(LIOB33_X0Y183_IOB_X0Y184_I),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_BO6),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f112f221f112f22)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_DLUT (
.I0(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f0000000)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_DLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800800080008000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_CLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af0f0f0a0000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000006ccccccc)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4080000000000000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_CLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I4(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6708060000000000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h808080806c6c6c6c)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe80000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AQ),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1e78871e80808080)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111ff112222ff22)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h366ccccc33366ccc)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8eff008e00000000)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa5af05af0)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6000000078006000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1fe07f8007f81fe0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2aa00a220aa0020)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I3(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.I5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a05a5a5a5a)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00ff00ff00)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5b7f32b3135b2032)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff00aa55aaaa55)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666699999999)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555c03f4015)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cccc33e0bbb0ee)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.I4(CLBLM_R_X11Y124_SLICE_X15Y124_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ddddffff)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.Q(CLBLM_R_X7Y107_SLICE_X8Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcf0cc00)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h030cabae030cabae)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0099f0f90066f0f6)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fffffa00fa)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00cfcc0f00cfcc)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66996699dd44dd44)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.I2(1'b1),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef00efefee00eeee)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33ff33ee22)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(LIOB33_X0Y147_IOB_X0Y148_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0008000a0000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff88ff88ff88)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcd3bffffcd09)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f030b0ffff33bb)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f300f300f3)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0fef6faf0fef6)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1fff1fffffff2f2)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff6996)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fbbaa0b0a)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefefefffcfcfc)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffafef0fc)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fff4fff4)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff0fff044)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I2(LIOB33_X0Y191_IOB_X0Y192_I),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa33ffaa00ee00)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbfbffffaafa)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f311f100300010)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0e0f0fc0e0ccee)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5f5f5f5)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff044fffff044)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff7f)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000be3c8200)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.Q(CLBLM_R_X7Y111_SLICE_X9Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeccaa00eeccaa00)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h053b221f3b051f22)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbabfbfbf303f3f3)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffccccff0a)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3303ff0f77777777)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff00ffff0f0f)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I1(1'b1),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000005050005)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0aff02ff)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa0aaa02aa)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfb0efa0a)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0e00440000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffb33fb33)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba3030ffbaff30)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaa0000f0ff)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_A5Q),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000700077)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fff4ffcfffcff)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccff000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000efff00001000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaa0aaccccffff)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdccccc00050000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfff000cc00f0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aa33aa33)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd55ddd555dd555dd)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5ea9d6eb976ab57)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb22bbbb2b22bb2b)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h23022302dcbddcfd)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffafffa0a0afa0a0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202080c02020206)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554545450505050)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(LIOB33_X0Y185_IOB_X0Y185_I),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0eeee)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe400e4fff000f0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ae00ffffaeae)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aae0eef0ffe0ee)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(CLBLM_R_X15Y107_SLICE_X21Y107_CQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfa0afa0a)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030303030)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf300f000f700f500)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.I2(LIOB33_X0Y185_IOB_X0Y185_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000408ffffaa55)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ffff4444)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff12ff)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000c004c4c4c4c)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003000001000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a2a2a2af5f5f5f5)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafa0000f0f0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff4f4f4fff444444)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff2f00000f2f0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.I3(LIOB33_X0Y161_IOB_X0Y161_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_B5Q),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb080baaaa0a0aaaa)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(LIOB33_X0Y165_IOB_X0Y165_I),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I5(LIOB33_X0Y185_IOB_X0Y185_I),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5ffd5c0c0ffc0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_B5Q),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff00cc80ffa0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(LIOB33_X0Y165_IOB_X0Y165_I),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbf00bfafaf00af)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I1(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aa66aa00000000)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbeefbfeaaaafafa)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffff008000a0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I2(LIOB33_X0Y157_IOB_X0Y158_I),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffaaccccfffa)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff030c030c030c)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3030ffffb8b8)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(LIOB33_X0Y159_IOB_X0Y160_I),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f41144f4f44444)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0f88880808)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5f5f5f5)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7373ffff4040)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(LIOB33_X0Y161_IOB_X0Y162_I),
.I3(1'b1),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5ffd5c0c0ffc0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0f88088808)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1230303030303030)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9333933380008000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h006c00cc005a00f0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa555580000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hae0cae0cae0cae0c)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3b3a0a0b3b3a0a0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(LIOB33_X0Y151_IOB_X0Y152_I),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf800f000f000f000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafa0afac)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(LIOB33_X0Y167_IOB_X0Y168_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0155015511551155)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffd500d5d5)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(LIOB33_X0Y159_IOB_X0Y159_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1115115511151155)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fdd0d5505)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0f22ff020f)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaafa00f000f0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(LIOB33_X0Y155_IOB_X0Y155_I),
.I1(1'b1),
.I2(LIOB33_X0Y171_IOB_X0Y171_I),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8ffc8ffc0ffc0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0fff0ccc8fffa)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(LIOB33_X0Y169_IOB_X0Y170_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011003300ff00ff)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcc0f00aa55aa55)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.I3(LIOB33_X0Y169_IOB_X0Y169_I),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ffdd0f050f0d)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a6a6a6a6a6a6a6a)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(LIOB33_X0Y169_IOB_X0Y170_I),
.I1(LIOB33_X0Y169_IOB_X0Y169_I),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h870f0f0f0f0f0f0f)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(LIOB33_X0Y171_IOB_X0Y172_I),
.I1(LIOB33_X0Y169_IOB_X0Y169_I),
.I2(LIOB33_X0Y173_IOB_X0Y173_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.I4(LIOB33_X0Y169_IOB_X0Y170_I),
.I5(LIOB33_X0Y171_IOB_X0Y171_I),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f066aaaaaa)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(LIOB33_X0Y171_IOB_X0Y171_I),
.I1(LIOB33_X0Y169_IOB_X0Y169_I),
.I2(LIOB33_X0Y171_IOB_X0Y172_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.I4(LIOB33_X0Y169_IOB_X0Y170_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f00ff0000000000)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.I1(LIOB33_X0Y177_IOB_X0Y178_I),
.I2(LIOB33_X0Y179_IOB_X0Y180_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(LIOB33_X0Y179_IOB_X0Y179_I),
.I5(LIOB33_X0Y181_IOB_X0Y181_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5f9f5f88008800)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(LIOB33_X0Y177_IOB_X0Y177_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(LIOB33_X0Y175_IOB_X0Y176_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cc0c0c048888888)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(LIOB33_X0Y179_IOB_X0Y180_I),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(LIOB33_X0Y179_IOB_X0Y179_I),
.I3(LIOB33_X0Y177_IOB_X0Y178_I),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb77bb770c0cc0c0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(LIOB33_X0Y177_IOB_X0Y178_I),
.I3(LIOB33_X0Y175_IOB_X0Y176_I),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h40c040c000000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.I1(LIOB33_X0Y173_IOB_X0Y174_I),
.I2(LIOB33_X0Y175_IOB_X0Y175_I),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y181_IOB_X0Y181_I),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d55f7ffdd5577ff)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(LIOB33_X0Y173_IOB_X0Y174_I),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.I3(LIOB33_X0Y181_IOB_X0Y181_I),
.I4(LIOB33_X0Y175_IOB_X0Y175_I),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3933333308000000)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(LIOB33_X0Y167_IOB_X0Y167_I),
.I1(LIOB33_X0Y167_IOB_X0Y168_I),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.I3(LIOB33_X0Y181_IOB_X0Y181_I),
.I4(LIOB33_X0Y165_IOB_X0Y166_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff8f8f033f)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(LIOB33_X0Y183_IOB_X0Y183_I),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf88ff0affffffff)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(LIOB33_X0Y185_IOB_X0Y185_I),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f351515151)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(LIOB33_X0Y173_IOB_X0Y173_I),
.I1(LIOB33_X0Y169_IOB_X0Y170_I),
.I2(1'b1),
.I3(LIOB33_X0Y171_IOB_X0Y172_I),
.I4(1'b1),
.I5(LIOB33_X0Y167_IOB_X0Y167_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000101)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(LIOB33_X0Y165_IOB_X0Y166_I),
.I1(LIOB33_X0Y169_IOB_X0Y169_I),
.I2(LIOB33_X0Y167_IOB_X0Y168_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_DO6),
.I5(LIOB33_X0Y171_IOB_X0Y171_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffc3ffc3ffc3ff)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y181_IOB_X0Y181_I),
.I2(LIOB33_X0Y173_IOB_X0Y174_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ccff3355995555)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(LIOB33_X0Y167_IOB_X0Y167_I),
.I1(LIOB33_X0Y181_IOB_X0Y181_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.I4(LIOB33_X0Y165_IOB_X0Y166_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y100_SLICE_X14Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y100_SLICE_X14Y100_DO5),
.O6(CLBLM_R_X11Y100_SLICE_X14Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_R_X11Y100_SLICE_X14Y100_CLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.O5(CLBLM_R_X11Y100_SLICE_X14Y100_CO5),
.O6(CLBLM_R_X11Y100_SLICE_X14Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y100_SLICE_X14Y100_BLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I5(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.O5(CLBLM_R_X11Y100_SLICE_X14Y100_BO5),
.O6(CLBLM_R_X11Y100_SLICE_X14Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f807f8080008000)
  ) CLBLM_R_X11Y100_SLICE_X14Y100_ALUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y100_SLICE_X14Y100_AO5),
.O6(CLBLM_R_X11Y100_SLICE_X14Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y100_SLICE_X15Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y100_SLICE_X15Y100_DO5),
.O6(CLBLM_R_X11Y100_SLICE_X15Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y100_SLICE_X15Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y100_SLICE_X15Y100_CO5),
.O6(CLBLM_R_X11Y100_SLICE_X15Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y100_SLICE_X15Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y100_SLICE_X15Y100_BO5),
.O6(CLBLM_R_X11Y100_SLICE_X15Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y100_SLICE_X15Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y100_SLICE_X15Y100_AO5),
.O6(CLBLM_R_X11Y100_SLICE_X15Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y101_SLICE_X14Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y101_SLICE_X14Y101_AO6),
.Q(CLBLM_R_X11Y101_SLICE_X14Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h56aa6aaaaaaaaaaa)
  ) CLBLM_R_X11Y101_SLICE_X14Y101_DLUT (
.I0(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I1(CLBLM_R_X11Y100_SLICE_X14Y100_AO5),
.I2(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I4(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.O5(CLBLM_R_X11Y101_SLICE_X14Y101_DO5),
.O6(CLBLM_R_X11Y101_SLICE_X14Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h055005503773cddc)
  ) CLBLM_R_X11Y101_SLICE_X14Y101_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_R_X11Y102_SLICE_X14Y102_AO5),
.I2(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I3(CLBLM_L_X10Y101_SLICE_X12Y101_AO6),
.I4(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_R_X11Y101_SLICE_X14Y101_CO5),
.O6(CLBLM_R_X11Y101_SLICE_X14Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000080000000)
  ) CLBLM_R_X11Y101_SLICE_X14Y101_BLUT (
.I0(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.O5(CLBLM_R_X11Y101_SLICE_X14Y101_BO5),
.O6(CLBLM_R_X11Y101_SLICE_X14Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffcfcf00cf)
  ) CLBLM_R_X11Y101_SLICE_X14Y101_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y101_SLICE_X15Y101_DO6),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I5(CLBLM_R_X11Y101_SLICE_X14Y101_CO6),
.O5(CLBLM_R_X11Y101_SLICE_X14Y101_AO5),
.O6(CLBLM_R_X11Y101_SLICE_X14Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3f0f3f0f3f0)
  ) CLBLM_R_X11Y101_SLICE_X15Y101_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I3(CLBLM_R_X11Y102_SLICE_X14Y102_AO5),
.I4(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X11Y101_SLICE_X15Y101_DO5),
.O6(CLBLM_R_X11Y101_SLICE_X15Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h003caabe00ccaaee)
  ) CLBLM_R_X11Y101_SLICE_X15Y101_CLUT (
.I0(CLBLM_R_X11Y101_SLICE_X15Y101_AO6),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_L_X10Y100_SLICE_X12Y100_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.O5(CLBLM_R_X11Y101_SLICE_X15Y101_CO5),
.O6(CLBLM_R_X11Y101_SLICE_X15Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y101_SLICE_X15Y101_BLUT (
.I0(CLBLM_R_X11Y100_SLICE_X14Y100_CO6),
.I1(CLBLM_R_X11Y102_SLICE_X14Y102_AO5),
.I2(CLBLM_R_X11Y100_SLICE_X14Y100_AO6),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.I4(CLBLM_R_X11Y101_SLICE_X15Y101_AO6),
.I5(CLBLM_R_X11Y101_SLICE_X15Y101_AO5),
.O5(CLBLM_R_X11Y101_SLICE_X15Y101_BO5),
.O6(CLBLM_R_X11Y101_SLICE_X15Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3fc03fc0)
  ) CLBLM_R_X11Y101_SLICE_X15Y101_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y101_SLICE_X15Y101_AO5),
.O6(CLBLM_R_X11Y101_SLICE_X15Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcceeccddccee)
  ) CLBLM_R_X11Y102_SLICE_X14Y102_DLUT (
.I0(CLBLM_L_X10Y100_SLICE_X12Y100_BO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X11Y102_SLICE_X14Y102_DO5),
.O6(CLBLM_R_X11Y102_SLICE_X14Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0affffff0a)
  ) CLBLM_R_X11Y102_SLICE_X14Y102_CLUT (
.I0(CLBLM_L_X12Y102_SLICE_X17Y102_AO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X11Y100_SLICE_X14Y100_CO6),
.I4(CLBLM_R_X11Y102_SLICE_X14Y102_DO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_R_X11Y102_SLICE_X14Y102_CO5),
.O6(CLBLM_R_X11Y102_SLICE_X14Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4080000000000000)
  ) CLBLM_R_X11Y102_SLICE_X14Y102_BLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I2(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.O5(CLBLM_R_X11Y102_SLICE_X14Y102_BO5),
.O6(CLBLM_R_X11Y102_SLICE_X14Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000078f0f0f0)
  ) CLBLM_R_X11Y102_SLICE_X14Y102_ALUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I2(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y102_SLICE_X14Y102_AO5),
.O6(CLBLM_R_X11Y102_SLICE_X14Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X11Y102_SLICE_X15Y102_DLUT (
.I0(CLBLM_L_X12Y102_SLICE_X17Y102_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y102_SLICE_X13Y102_CO6),
.O5(CLBLM_R_X11Y102_SLICE_X15Y102_DO5),
.O6(CLBLM_R_X11Y102_SLICE_X15Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b0a3b0a3b0a3b0a)
  ) CLBLM_R_X11Y102_SLICE_X15Y102_CLUT (
.I0(CLBLM_R_X11Y102_SLICE_X15Y102_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X11Y103_SLICE_X15Y103_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y102_SLICE_X15Y102_CO5),
.O6(CLBLM_R_X11Y102_SLICE_X15Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y102_SLICE_X15Y102_BLUT (
.I0(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I1(CLBLM_L_X12Y102_SLICE_X17Y102_AO6),
.I2(CLBLM_L_X10Y103_SLICE_X13Y103_AO6),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I4(CLBLM_R_X11Y102_SLICE_X15Y102_AO6),
.I5(CLBLM_R_X11Y102_SLICE_X15Y102_AO5),
.O5(CLBLM_R_X11Y102_SLICE_X15Y102_BO5),
.O6(CLBLM_R_X11Y102_SLICE_X15Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cccccc55aaff00)
  ) CLBLM_R_X11Y102_SLICE_X15Y102_ALUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I1(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y102_SLICE_X15Y102_AO5),
.O6(CLBLM_R_X11Y102_SLICE_X15Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y103_SLICE_X14Y103_AO6),
.Q(CLBLM_R_X11Y103_SLICE_X14Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdedededeedededed)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_DLUT (
.I0(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_DO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf232300000000)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I2(CLBLM_R_X11Y103_SLICE_X15Y103_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(CLBLM_R_X11Y103_SLICE_X14Y103_DO6),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_CO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000099090000)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_BLUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I1(CLBLM_R_X11Y102_SLICE_X14Y102_AO5),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_BO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h75ff000075ff75ff)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_ALUT (
.I0(CLBLM_R_X11Y103_SLICE_X14Y103_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I2(CLBLM_R_X11Y103_SLICE_X15Y103_DO6),
.I3(CLBLM_R_X11Y103_SLICE_X14Y103_BO6),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_AO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa5555aaaa)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_DLUT (
.I0(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_DO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f030f0305010501)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_CLUT (
.I0(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I1(CLBLM_R_X11Y102_SLICE_X15Y102_DO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_CO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1fe07f80ff00ff00)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_BLUT (
.I0(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I4(CLBLM_R_X11Y101_SLICE_X14Y101_AQ),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_BO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cca5ed5ade)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_ALUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I1(CLBLM_R_X11Y102_SLICE_X15Y102_DO6),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_AO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.Q(CLBLM_R_X11Y104_SLICE_X14Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa000fffa0000)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_DLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffb3a0)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AQ),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbabaffba)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffe0f0a0f0e)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_BO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cc0c0000ff0f)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_R_X11Y103_SLICE_X15Y103_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I4(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcecffffdcecdcec)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f228f88afaa0f00)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f80ff00ff00ff00)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I3(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I4(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I3(CLBLM_L_X12Y103_SLICE_X16Y103_AQ),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ba30baba30ba30)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000022)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000100)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00ff91)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y103_SLICE_X11Y103_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f066666666)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefafffffeeaa)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaff0000283c)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff2f11)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaaba)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0f0f2)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5055055510110111)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00033ccff00)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_AQ),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffceffffcece)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffeeffcfffcc)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I1(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I5(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080a0aa88)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafefaabb)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33b733b700a500a5)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h001e000f00660033)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfb00fbfbfb00fb)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I1(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ffbb0f030f0b)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffc0003fff)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5577003377553300)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000000a)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff95555555)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf8a454545)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22112211cfcffcfc)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ffc0cc3033)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000055a500003363)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f351f3f3f351)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y195_IOB_X0Y195_I),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h007f0080007f0080)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_CLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcced0021ffff3333)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y112_SLICE_X15Y112_AO6),
.Q(CLBLM_R_X11Y112_SLICE_X15Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_DLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_CLUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000080000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_BLUT (
.I0(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff0033deff1233)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000000000000)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h35ff70ff35357070)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc0080808080)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I1(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaa03030303)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafbbbfaa0f333f00)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_A5Q),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000055aa000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I3(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I4(CLBLM_L_X12Y114_SLICE_X17Y114_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h507350dcdcffdcdc)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcddc0550ffdcff50)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_A5Q),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_A5Q),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I5(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afcfc0c0c)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_AO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.Q(CLBLM_R_X11Y114_SLICE_X15Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeedddd00ee00dd)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f7f33775f0f5500)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff78)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_A5Q),
.I2(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_DO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff00080808080)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fcfcf0000cccc)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50507c7cff50ff7c)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaa12aa30)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f11dfdd4f44cfcc)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I2(CLBLM_R_X11Y124_SLICE_X15Y124_AO6),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I3(CLBLM_R_X11Y114_SLICE_X15Y114_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_A5Q),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffaaff0000aaaa)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heefcaa30eefcaa30)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88f3f3c0c0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_A5Q),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f8f8f8f88888888)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BQ),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1122f1f2bbaafbfa)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_A5Q),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f300f077f7aafa)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.I4(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55aa00be50)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_CO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffe)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ace0a0aff3b0a0a)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c5d5d0cffff5d0c)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f4f4fff4444ff44)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_A5Q),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(LIOB33_X0Y147_IOB_X0Y147_I),
.I1(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_BO6),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fcfcfff0fffc)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0a44444e4e)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa2222faaa3222)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y151_IOB_X0Y151_I),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_BO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_CO6),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff00fffcfff0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000001)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aaa0aae0eea0aa)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888f8f8f8f8)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.I2(LIOB33_X0Y155_IOB_X0Y155_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff44fff4fff4)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b3f5f5a0b3a0a0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ff08080008)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(LIOB33_X0Y151_IOB_X0Y152_I),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_CO6),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0cff0fdddddddd)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b038bcfcc00cc00)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330033f0bbf088)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(CLBLM_R_X13Y124_SLICE_X18Y124_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_L_X12Y125_SLICE_X17Y125_BO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X13Y120_SLICE_X18Y120_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddf5a08888f5a0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_BO6),
.I3(CLBLM_R_X13Y120_SLICE_X19Y120_BO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb051105bbaf11af)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_R_X13Y120_SLICE_X19Y120_DO6),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa30fa3f0a300a3)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X19Y120_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.I5(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa303f0a0a303f)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(CLBLM_R_X13Y120_SLICE_X19Y120_DO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaf0faf0fa)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h333333330055aaff)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_CO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_BO6),
.I4(CLBLM_L_X12Y124_SLICE_X16Y124_DO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbf3bbc088f388c0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_R_X13Y120_SLICE_X19Y120_DO6),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0f550fff0000ff)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_DO6),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_CO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaabbaa33003300)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_BO5),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y157_IOB_X0Y157_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_CO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacfff0acac0f00)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_DO6),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X12Y125_SLICE_X17Y125_AO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X17Y125_AO6),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcff505c0c0f505)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(CLBLM_R_X13Y124_SLICE_X18Y124_DO6),
.I1(CLBLM_L_X12Y125_SLICE_X17Y125_AO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y120_SLICE_X18Y120_DO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ff55550f0f)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05af058888dddd)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccfff0aacc00f0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_CO6),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.I2(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaf0caffca00ca0f)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfafc0a0cfa0c0a)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0434c4f40737c7f7)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.I4(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_CO6),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30503f50305f3f5f)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(CLBLM_L_X12Y123_SLICE_X16Y123_AQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fafaee445050)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_L_X12Y124_SLICE_X16Y124_CO6),
.I2(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5ee44a0a0ee44)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_CO6),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0c5c50f00c5c5)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_DO6),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X13Y121_SLICE_X18Y121_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X13Y125_SLICE_X19Y125_BO6),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33fd31fc30)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_CO6),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I4(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff40ffff404040)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I4(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffeaeac0ff)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000010000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffaaccccfffa)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.I1(CLBLM_R_X15Y120_SLICE_X21Y120_AQ),
.I2(LIOB33_X0Y157_IOB_X0Y157_I),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_DO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10b01aba15b51fbf)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X16Y126_SLICE_X22Y126_AQ),
.I4(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff0facacf000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I1(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_L_X16Y126_SLICE_X22Y126_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200100000)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa003300aaff33ff)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeaa44554400)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_L_X12Y124_SLICE_X17Y124_CO6),
.I5(CLBLM_R_X11Y124_SLICE_X15Y124_BO6),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h11110111ddddcddd)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0f3f3afa00303)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_DO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_L_X12Y124_SLICE_X17Y124_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5353535300f00fff)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I1(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffb1b1ffb1)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(LIOB33_X0Y153_IOB_X0Y153_I),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_CO6),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afe0efe0e)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y125_SLICE_X15Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X15Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ddddfa508888)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03cf03cf03cf02ce)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_R_X13Y125_SLICE_X19Y125_DO6),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0f3c0fbea)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I2(CLBLM_R_X11Y125_SLICE_X15Y125_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff0fffa)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_BO6),
.I3(CLBLM_R_X11Y125_SLICE_X15Y125_BO6),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffddccffff5f0f)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_CLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_DO6),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033ff3b0a3b)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555bbaa1100)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_CO6),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffaaf0cc00aaf0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_DLUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3355000f3355ff0f)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_CLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I2(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h05af05af1111bbbb)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0eff0ffe0efe0e)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X12Y126_SLICE_X17Y126_AQ),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I5(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_BO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bb00bb0b0b0b0b)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_BQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0555055503330333)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I4(1'b1),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1f3d1d1f3f3f3f3)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X14Y127_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1f3d1d1f3f3f3f3)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefc302222fc30)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_DLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c3f11110c3fdddd)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_CLUT (
.I0(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000080000)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000001)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55cc55ccffff55cc)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I4(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff04ffffff02ff)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_BO6),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000004fffbffff)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffae00ff00ae)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.I1(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I2(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c008c00af23af23)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I2(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h40400000fffffffd)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000010ffffefff)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfdffff11313333)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y153_IOB_X0Y153_I),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.I5(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3bbf388c0bbc088)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_DLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0311cf1103ddcfdd)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_CLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b3f5f7a0a0f5f5)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffddf0f0ffcc)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.I2(CLBLM_L_X12Y124_SLICE_X16Y124_AQ),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y129_SLICE_X15Y129_BO6),
.Q(CLBLM_R_X11Y129_SLICE_X15Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeaadd55cc00)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_DLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I4(CLBLM_R_X11Y129_SLICE_X15Y129_AQ),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77335500ffbbffaa)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_CLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_BQ),
.I4(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffba5510)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_CO6),
.I2(LIOB33_X0Y151_IOB_X0Y152_I),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_AQ),
.I5(CLBLM_R_X11Y129_SLICE_X15Y129_CO6),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0aaf0fff0ee)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_ALUT (
.I0(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y129_SLICE_X21Y129_AO5),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_DO6),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbaaa3000baaa)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_AQ),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfefcfecceeffff)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_DO6),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_BO6),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88ddd8ddd8)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y125_SLICE_X16Y125_BQ),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_BO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y130_SLICE_X15Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X15Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3f0f33003f0f)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_AQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfaf3705)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I5(CLBLM_R_X11Y130_SLICE_X15Y130_CO6),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333efee2322)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_CO6),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffb00000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcccdcccd)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff5fd)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffe55445554)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_CO6),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_BO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I5(LIOB33_X0Y143_IOB_X0Y143_I),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3bfa0afb3bfa0af)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3e2e2e2f3)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ddd8ddd8)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(LIOB33_X0Y189_IOB_X0Y189_I),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_BO6),
.I3(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I4(1'b1),
.I5(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y100_SLICE_X18Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y100_SLICE_X18Y100_AO6),
.Q(CLBLM_R_X13Y100_SLICE_X18Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fcc330c03)
  ) CLBLM_R_X13Y100_SLICE_X18Y100_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I2(CLBLM_R_X13Y100_SLICE_X19Y100_BO6),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_CO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_R_X13Y100_SLICE_X18Y100_DO5),
.O6(CLBLM_R_X13Y100_SLICE_X18Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y100_SLICE_X18Y100_CLUT (
.I0(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I1(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I2(CLBLM_L_X10Y100_SLICE_X12Y100_BO6),
.I3(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.O5(CLBLM_R_X13Y100_SLICE_X18Y100_CO5),
.O6(CLBLM_R_X13Y100_SLICE_X18Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f088ccaaff)
  ) CLBLM_R_X13Y100_SLICE_X18Y100_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I2(CLBLM_L_X12Y101_SLICE_X17Y101_CO6),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_BO6),
.I4(CLBLM_R_X15Y100_SLICE_X20Y100_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y100_SLICE_X18Y100_BO5),
.O6(CLBLM_R_X13Y100_SLICE_X18Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd8ddd8ddd)
  ) CLBLM_R_X13Y100_SLICE_X18Y100_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_BO5),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_DO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y104_SLICE_X18Y104_CO6),
.O5(CLBLM_R_X13Y100_SLICE_X18Y100_AO5),
.O6(CLBLM_R_X13Y100_SLICE_X18Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y100_SLICE_X19Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y100_SLICE_X19Y100_DO5),
.O6(CLBLM_R_X13Y100_SLICE_X19Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y100_SLICE_X19Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y100_SLICE_X19Y100_CO5),
.O6(CLBLM_R_X13Y100_SLICE_X19Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaaaaaaaaaaaaaa)
  ) CLBLM_R_X13Y100_SLICE_X19Y100_BLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I2(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I3(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I5(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.O5(CLBLM_R_X13Y100_SLICE_X19Y100_BO5),
.O6(CLBLM_R_X13Y100_SLICE_X19Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y100_SLICE_X19Y100_ALUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I2(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I4(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I5(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.O5(CLBLM_R_X13Y100_SLICE_X19Y100_AO5),
.O6(CLBLM_R_X13Y100_SLICE_X19Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y101_SLICE_X18Y101_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y101_SLICE_X18Y101_AO6),
.Q(CLBLM_R_X13Y101_SLICE_X18Y101_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cff0cff0c0c0c0c)
  ) CLBLM_R_X13Y101_SLICE_X18Y101_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y101_SLICE_X19Y101_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y102_SLICE_X17Y102_BO6),
.O5(CLBLM_R_X13Y101_SLICE_X18Y101_DO5),
.O6(CLBLM_R_X13Y101_SLICE_X18Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a3b0ace0a3b0ace)
  ) CLBLM_R_X13Y101_SLICE_X18Y101_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X19Y102_AO6),
.I1(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_R_X13Y101_SLICE_X18Y101_BO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y101_SLICE_X18Y101_CO5),
.O6(CLBLM_R_X13Y101_SLICE_X18Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X13Y101_SLICE_X18Y101_BLUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I2(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I3(CLBLM_L_X10Y100_SLICE_X12Y100_BO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y101_SLICE_X18Y101_BO5),
.O6(CLBLM_R_X13Y101_SLICE_X18Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff0eef0ee)
  ) CLBLM_R_X13Y101_SLICE_X18Y101_ALUT (
.I0(CLBLM_R_X13Y103_SLICE_X18Y103_DO6),
.I1(CLBLM_R_X13Y101_SLICE_X18Y101_DO6),
.I2(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y101_SLICE_X18Y101_CO6),
.O5(CLBLM_R_X13Y101_SLICE_X18Y101_AO5),
.O6(CLBLM_R_X13Y101_SLICE_X18Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y101_SLICE_X19Y101_DLUT (
.I0(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I1(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I3(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I4(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I5(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.O5(CLBLM_R_X13Y101_SLICE_X19Y101_DO5),
.O6(CLBLM_R_X13Y101_SLICE_X19Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y101_SLICE_X19Y101_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X19Y102_AO6),
.I1(CLBLM_R_X13Y100_SLICE_X19Y100_BO6),
.I2(CLBLM_R_X13Y103_SLICE_X19Y103_AO6),
.I3(CLBLM_R_X15Y101_SLICE_X21Y101_BO5),
.I4(CLBLM_R_X15Y101_SLICE_X20Y101_AO5),
.I5(CLBLM_R_X11Y101_SLICE_X15Y101_BO6),
.O5(CLBLM_R_X13Y101_SLICE_X19Y101_CO5),
.O6(CLBLM_R_X13Y101_SLICE_X19Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y101_SLICE_X19Y101_BLUT (
.I0(CLBLM_R_X15Y101_SLICE_X21Y101_AO5),
.I1(CLBLM_R_X11Y102_SLICE_X15Y102_BO6),
.I2(CLBLM_R_X15Y100_SLICE_X20Y100_BO6),
.I3(CLBLM_R_X15Y101_SLICE_X20Y101_BO5),
.I4(CLBLM_R_X13Y101_SLICE_X19Y101_AO6),
.I5(CLBLM_R_X13Y103_SLICE_X19Y103_CO6),
.O5(CLBLM_R_X13Y101_SLICE_X19Y101_BO5),
.O6(CLBLM_R_X13Y101_SLICE_X19Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff800080000000)
  ) CLBLM_R_X13Y101_SLICE_X19Y101_ALUT (
.I0(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I2(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I3(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I4(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y101_SLICE_X19Y101_AO5),
.O6(CLBLM_R_X13Y101_SLICE_X19Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y102_SLICE_X18Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y102_SLICE_X18Y102_AO6),
.Q(CLBLM_R_X13Y102_SLICE_X18Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X13Y102_SLICE_X18Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y102_SLICE_X17Y102_DO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y103_SLICE_X19Y103_AO6),
.O5(CLBLM_R_X13Y102_SLICE_X18Y102_DO5),
.O6(CLBLM_R_X13Y102_SLICE_X18Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f3f0fcf003300cc)
  ) CLBLM_R_X13Y102_SLICE_X18Y102_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y103_SLICE_X17Y103_CO6),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLM_R_X13Y103_SLICE_X19Y103_CO6),
.I5(CLBLM_R_X13Y103_SLICE_X19Y103_AO6),
.O5(CLBLM_R_X13Y102_SLICE_X18Y102_CO5),
.O6(CLBLM_R_X13Y102_SLICE_X18Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3311331130100301)
  ) CLBLM_R_X13Y102_SLICE_X18Y102_BLUT (
.I0(CLBLM_R_X13Y103_SLICE_X19Y103_CO6),
.I1(CLBLM_R_X13Y103_SLICE_X18Y103_BO6),
.I2(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLM_R_X13Y101_SLICE_X18Y101_BO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_R_X13Y102_SLICE_X18Y102_BO5),
.O6(CLBLM_R_X13Y102_SLICE_X18Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0ff55555055)
  ) CLBLM_R_X13Y102_SLICE_X18Y102_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(1'b1),
.I2(CLBLM_R_X13Y103_SLICE_X19Y103_DO6),
.I3(CLBLM_R_X13Y102_SLICE_X18Y102_BO6),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_CO6),
.I5(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.O5(CLBLM_R_X13Y102_SLICE_X18Y102_AO5),
.O6(CLBLM_R_X13Y102_SLICE_X18Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff09ff06ff09ff06)
  ) CLBLM_R_X13Y102_SLICE_X19Y102_DLUT (
.I0(CLBLM_R_X15Y102_SLICE_X21Y102_AO6),
.I1(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_R_X13Y102_SLICE_X19Y102_CO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y102_SLICE_X19Y102_DO5),
.O6(CLBLM_R_X13Y102_SLICE_X19Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000001f7fe080)
  ) CLBLM_R_X13Y102_SLICE_X19Y102_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_L_X12Y102_SLICE_X17Y102_DO6),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X13Y102_SLICE_X19Y102_AO5),
.I4(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.O5(CLBLM_R_X13Y102_SLICE_X19Y102_CO5),
.O6(CLBLM_R_X13Y102_SLICE_X19Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77887f807f80ff00)
  ) CLBLM_R_X13Y102_SLICE_X19Y102_BLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I2(CLBLM_L_X12Y102_SLICE_X17Y102_DO6),
.I3(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I5(CLBLM_R_X13Y102_SLICE_X19Y102_AO5),
.O5(CLBLM_R_X13Y102_SLICE_X19Y102_BO5),
.O6(CLBLM_R_X13Y102_SLICE_X19Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccccccc0000000)
  ) CLBLM_R_X13Y102_SLICE_X19Y102_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I2(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I3(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y102_SLICE_X19Y102_AO5),
.O6(CLBLM_R_X13Y102_SLICE_X19Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y103_SLICE_X18Y103_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y103_SLICE_X18Y103_AO6),
.Q(CLBLM_R_X13Y103_SLICE_X18Y103_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffb3a0)
  ) CLBLM_R_X13Y103_SLICE_X18Y103_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I3(CLBLM_L_X12Y102_SLICE_X17Y102_CO6),
.I4(CLBLM_R_X15Y108_SLICE_X20Y108_CO6),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_DO6),
.O5(CLBLM_R_X13Y103_SLICE_X18Y103_DO5),
.O6(CLBLM_R_X13Y103_SLICE_X18Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfafffffbbaa)
  ) CLBLM_R_X13Y103_SLICE_X18Y103_CLUT (
.I0(CLBLM_R_X13Y107_SLICE_X18Y107_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I3(CLBLM_L_X12Y102_SLICE_X17Y102_CO6),
.I4(CLBLM_R_X15Y108_SLICE_X20Y108_CO6),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.O5(CLBLM_R_X13Y103_SLICE_X18Y103_CO5),
.O6(CLBLM_R_X13Y103_SLICE_X18Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3003033021222212)
  ) CLBLM_R_X13Y103_SLICE_X18Y103_BLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_L_X12Y103_SLICE_X17Y103_BO6),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y103_SLICE_X18Y103_BO5),
.O6(CLBLM_R_X13Y103_SLICE_X18Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf070ff77f030ff33)
  ) CLBLM_R_X13Y103_SLICE_X18Y103_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I1(CLBLM_R_X13Y103_SLICE_X19Y103_BO6),
.I2(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I3(CLBLM_R_X13Y103_SLICE_X18Y103_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y102_SLICE_X18Y102_DO6),
.O5(CLBLM_R_X13Y103_SLICE_X18Y103_AO5),
.O6(CLBLM_R_X13Y103_SLICE_X18Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaeeffff00cc)
  ) CLBLM_R_X13Y103_SLICE_X19Y103_DLUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_R_X13Y102_SLICE_X18Y102_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_R_X15Y108_SLICE_X20Y108_BO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X13Y103_SLICE_X19Y103_DO5),
.O6(CLBLM_R_X13Y103_SLICE_X19Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaaaaaaaaaaaaaa)
  ) CLBLM_R_X13Y103_SLICE_X19Y103_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I4(CLBLM_L_X12Y102_SLICE_X16Y102_AQ),
.I5(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.O5(CLBLM_R_X13Y103_SLICE_X19Y103_CO5),
.O6(CLBLM_R_X13Y103_SLICE_X19Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a080f0c080a0c0f)
  ) CLBLM_R_X13Y103_SLICE_X19Y103_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I2(CLBLM_R_X13Y106_SLICE_X19Y106_AO6),
.I3(CLBLM_L_X12Y103_SLICE_X17Y103_CO6),
.I4(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I5(CLBLM_R_X13Y103_SLICE_X19Y103_CO6),
.O5(CLBLM_R_X13Y103_SLICE_X19Y103_BO5),
.O6(CLBLM_R_X13Y103_SLICE_X19Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f080000000)
  ) CLBLM_R_X13Y103_SLICE_X19Y103_ALUT (
.I0(CLBLM_L_X12Y101_SLICE_X16Y101_BQ),
.I1(CLBLM_L_X12Y102_SLICE_X16Y102_BQ),
.I2(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I3(CLBLM_R_X11Y100_SLICE_X14Y100_BO6),
.I4(CLBLM_R_X13Y101_SLICE_X18Y101_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y103_SLICE_X19Y103_AO5),
.O6(CLBLM_R_X13Y103_SLICE_X19Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y104_SLICE_X18Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y104_SLICE_X18Y104_AO6),
.Q(CLBLM_R_X13Y104_SLICE_X18Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X13Y104_SLICE_X18Y104_DLUT (
.I0(CLBLM_L_X12Y101_SLICE_X17Y101_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X13Y100_SLICE_X19Y100_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y104_SLICE_X18Y104_DO5),
.O6(CLBLM_R_X13Y104_SLICE_X18Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffb3ffa0)
  ) CLBLM_R_X13Y104_SLICE_X18Y104_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X13Y103_SLICE_X18Y103_BO5),
.I4(CLBLM_R_X13Y104_SLICE_X18Y104_DO6),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_DO6),
.O5(CLBLM_R_X13Y104_SLICE_X18Y104_CO5),
.O6(CLBLM_R_X13Y104_SLICE_X18Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffeefffcfffe)
  ) CLBLM_R_X13Y104_SLICE_X18Y104_BLUT (
.I0(CLBLM_R_X13Y104_SLICE_X18Y104_DO6),
.I1(CLBLM_R_X13Y106_SLICE_X18Y106_DO6),
.I2(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_R_X13Y104_SLICE_X18Y104_BO5),
.O6(CLBLM_R_X13Y104_SLICE_X18Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5a0f5e4)
  ) CLBLM_R_X13Y104_SLICE_X18Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y100_SLICE_X18Y100_BO6),
.I2(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I3(CLBLM_R_X13Y104_SLICE_X18Y104_BO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(CLBLM_R_X13Y103_SLICE_X18Y103_BO5),
.O5(CLBLM_R_X13Y104_SLICE_X18Y104_AO5),
.O6(CLBLM_R_X13Y104_SLICE_X18Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y104_SLICE_X19Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y104_SLICE_X19Y104_AO6),
.Q(CLBLM_R_X13Y104_SLICE_X19Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y104_SLICE_X19Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y104_SLICE_X19Y104_DO5),
.O6(CLBLM_R_X13Y104_SLICE_X19Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y104_SLICE_X19Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y104_SLICE_X19Y104_CO5),
.O6(CLBLM_R_X13Y104_SLICE_X19Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y104_SLICE_X19Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y104_SLICE_X19Y104_BO5),
.O6(CLBLM_R_X13Y104_SLICE_X19Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0faaee0a0e)
  ) CLBLM_R_X13Y104_SLICE_X19Y104_ALUT (
.I0(CLBLM_R_X13Y102_SLICE_X19Y102_DO6),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I4(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I5(CLBLM_R_X13Y106_SLICE_X18Y106_CO6),
.O5(CLBLM_R_X13Y104_SLICE_X19Y104_AO5),
.O6(CLBLM_R_X13Y104_SLICE_X19Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0cffc0000cccc)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y107_SLICE_X18Y107_BO6),
.I2(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I3(CLBLM_R_X13Y106_SLICE_X18Y106_AO5),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_DO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00f0ccfc)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y109_SLICE_X19Y109_AO6),
.I2(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(CLBLM_R_X13Y106_SLICE_X18Y106_BO6),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_CO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeffeaff0cffc0)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X13Y106_SLICE_X18Y106_AO6),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_BO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_ALUT (
.I0(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I2(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I4(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_AO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_DO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_CO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_BO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f5fdf5f3f0fcf0)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_AO6),
.I2(CLBLM_R_X15Y108_SLICE_X20Y108_BO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I5(CLBLM_R_X13Y107_SLICE_X18Y107_AO5),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_AO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cbe00aaf0fa00aa)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_DLUT (
.I0(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I2(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_DO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_CLUT (
.I0(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I1(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I3(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I4(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_CO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaaaaaaaaaaaaaa)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_BLUT (
.I0(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I2(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I4(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I5(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_BO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7f80807f80ff00)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_ALUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_AQ),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I2(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I3(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I4(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_AO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_DO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_CO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_BO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_AO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.Q(CLBLM_R_X13Y108_SLICE_X18Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000100)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_CLUT (
.I0(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I2(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I4(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000010)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_BLUT (
.I0(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I1(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.I4(CLBLM_L_X12Y104_SLICE_X16Y104_BQ),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454fefe5454)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_BO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5d5d5c0c0c0c0)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_DLUT (
.I0(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(CLBLM_R_X13Y104_SLICE_X18Y104_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X13Y107_SLICE_X18Y107_BO6),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4f44ffff444f)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I2(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I3(CLBLM_R_X13Y108_SLICE_X19Y108_AO5),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_DO6),
.I5(CLBLM_R_X13Y107_SLICE_X18Y107_BO6),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00f0ffff99f9)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_BLUT (
.I0(CLBLM_R_X13Y107_SLICE_X18Y107_AO5),
.I1(CLBLM_R_X13Y109_SLICE_X19Y109_BO6),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_AO6),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2222255005500)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_ALUT (
.I0(CLBLM_R_X13Y107_SLICE_X18Y107_AO5),
.I1(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(CLBLM_R_X13Y109_SLICE_X19Y109_BO6),
.I4(CLBLM_R_X13Y103_SLICE_X18Y103_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022222222)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_CLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I1(CLBLM_R_X13Y109_SLICE_X19Y109_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y108_SLICE_X20Y108_AO5),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00ccf0fc0fcf)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_AO6),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h444444444ff444ff)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_AO6),
.I3(CLBLM_R_X15Y108_SLICE_X20Y108_AO5),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I5(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0c0c0c0c)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_DO6),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y110_SLICE_X18Y110_AO6),
.Q(CLBLM_R_X13Y110_SLICE_X18Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffceffffff0a)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_DLUT (
.I0(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_AQ),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5d0cffff0c5d)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_CLUT (
.I0(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I1(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(CLBLM_L_X16Y109_SLICE_X23Y109_AO5),
.I4(CLBLM_R_X13Y112_SLICE_X18Y112_BO5),
.I5(CLBLM_R_X15Y110_SLICE_X21Y110_DO6),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbaabfafb)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_BLUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_DO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_DO6),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(CLBLM_L_X12Y112_SLICE_X17Y112_AO6),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ffd0ddd0dd)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_ALUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_DO6),
.I1(CLBLM_R_X15Y110_SLICE_X20Y110_DO6),
.I2(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y110_SLICE_X18Y110_CO6),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y111_SLICE_X18Y111_AO6),
.Q(CLBLM_R_X13Y111_SLICE_X18Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_DO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_CLUT (
.I0(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_CO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h02000000fffbfffb)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I4(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffce3302ffff3333)
  ) CLBLM_R_X13Y111_SLICE_X18Y111_ALUT (
.I0(CLBLM_R_X13Y109_SLICE_X19Y109_AO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_BO6),
.I4(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I5(CLBLM_R_X13Y114_SLICE_X18Y114_BO6),
.O5(CLBLM_R_X13Y111_SLICE_X18Y111_AO5),
.O6(CLBLM_R_X13Y111_SLICE_X18Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_DO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800000000000)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_CLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.I2(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_CO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd0d0d0d0dddd)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I3(1'b1),
.I4(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_CO6),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_BO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X13Y111_SLICE_X19Y111_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I2(CLBLM_L_X16Y109_SLICE_X22Y109_DO6),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X13Y111_SLICE_X19Y111_AO5),
.O6(CLBLM_R_X13Y111_SLICE_X19Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaff82c382c3)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I1(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I2(CLBLM_R_X15Y112_SLICE_X20Y112_AO5),
.I3(CLBLM_L_X12Y115_SLICE_X16Y115_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff10ff23)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_CLUT (
.I0(CLBLM_L_X16Y109_SLICE_X23Y109_AO5),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_R_X15Y110_SLICE_X21Y110_DO6),
.I3(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.I4(CLBLM_L_X16Y109_SLICE_X22Y109_DO6),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_BO6),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1023102321212121)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_BLUT (
.I0(CLBLM_L_X12Y115_SLICE_X16Y115_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I2(CLBLM_R_X13Y112_SLICE_X19Y112_CO6),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030000300200000)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_ALUT (
.I0(CLBLM_R_X15Y107_SLICE_X21Y107_CQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000004)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_CLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_CO6),
.I2(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I3(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033013200330033)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I4(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.I5(CLBLM_R_X13Y115_SLICE_X18Y115_CO6),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_ALUT (
.I0(CLBLM_L_X16Y109_SLICE_X22Y109_DO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y113_SLICE_X18Y113_AO6),
.Q(CLBLM_R_X13Y113_SLICE_X18Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y113_SLICE_X18Y113_BO6),
.Q(CLBLM_R_X13Y113_SLICE_X18Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa8222ffffc333)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I2(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa802affffc03f)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I1(CLBLM_R_X15Y112_SLICE_X20Y112_AO5),
.I2(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_AQ),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0fcaaaaffff)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_BLUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(CLBLM_R_X13Y112_SLICE_X18Y112_CO6),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y113_SLICE_X18Y113_CO6),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fffdd0f0d)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_ALUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_DO6),
.I1(CLBLM_R_X15Y110_SLICE_X20Y110_CO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X13Y114_SLICE_X18Y114_AO6),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I5(CLBLM_R_X13Y109_SLICE_X18Y109_AO6),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y113_SLICE_X19Y113_AO6),
.Q(CLBLM_R_X13Y113_SLICE_X19Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff887700ff)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_DLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.I2(1'b1),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000008afc0000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I2(CLBLM_R_X13Y114_SLICE_X18Y114_AO5),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I4(CLBLM_R_X13Y113_SLICE_X19Y113_DO6),
.I5(CLBLM_R_X15Y110_SLICE_X20Y110_AO6),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f53131f000f000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_BO6),
.I4(CLBLM_L_X12Y113_SLICE_X17Y113_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccffccf54455445)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I2(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.I3(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_DO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050000)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_CO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00a000a200a8)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_BLUT (
.I0(CLBLM_R_X13Y114_SLICE_X18Y114_DO6),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_BO6),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_BO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000004fb00040004)
  ) CLBLM_R_X13Y114_SLICE_X18Y114_ALUT (
.I0(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X18Y114_AO5),
.O6(CLBLM_R_X13Y114_SLICE_X18Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y114_SLICE_X19Y114_AO6),
.Q(CLBLM_R_X13Y114_SLICE_X19Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_DO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_CO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffcfcfffcff)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_BO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b0bbbbaa00aa00)
  ) CLBLM_R_X13Y114_SLICE_X19Y114_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I3(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y114_SLICE_X19Y114_AO5),
.O6(CLBLM_R_X13Y114_SLICE_X19Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y115_SLICE_X18Y115_AO6),
.Q(CLBLM_R_X13Y115_SLICE_X18Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ccccccccccccccc)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_DLUT (
.I0(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I1(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_DO6),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_DO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_CLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I2(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_A5Q),
.I4(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I5(CLBLM_L_X12Y116_SLICE_X17Y116_BQ),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_CO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f00bfaa0f33afbb)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_BLUT (
.I0(CLBLM_R_X13Y115_SLICE_X18Y115_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I3(CLBLM_L_X12Y116_SLICE_X16Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_BO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff088888888)
  ) CLBLM_R_X13Y115_SLICE_X18Y115_ALUT (
.I0(CLBLM_L_X16Y115_SLICE_X22Y115_BO6),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I2(CLBLM_R_X13Y108_SLICE_X19Y108_CO6),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X18Y115_AO5),
.O6(CLBLM_R_X13Y115_SLICE_X18Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_DO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_CO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_BO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y115_SLICE_X19Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y115_SLICE_X19Y115_AO5),
.O6(CLBLM_R_X13Y115_SLICE_X19Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y117_SLICE_X18Y117_AO6),
.Q(CLBLM_R_X13Y117_SLICE_X18Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3d1f3d1f3c0)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_ALUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y195_IOB_X0Y196_I),
.I3(CLBLM_L_X16Y117_SLICE_X23Y117_BO6),
.I4(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I5(CLBLM_R_X13Y115_SLICE_X18Y115_AO5),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0000f000000f00)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_AO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfefeffccffee)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_DLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_DO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_CLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_CO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000505f5f5ffff)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffc8fa88aa)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_ALUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_DO6),
.I1(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_CO6),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_AO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_DO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_CO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_BO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_AO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y120_SLICE_X18Y120_AO6),
.Q(CLBLM_R_X13Y120_SLICE_X18Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h353500f035350fff)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_DLUT (
.I0(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I1(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X15Y120_SLICE_X20Y120_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_L_X16Y121_SLICE_X22Y121_AQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3c0fffffbea)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_CLUT (
.I0(LIOB33_X0Y155_IOB_X0Y155_I),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebadc9876325410)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLM_R_X13Y120_SLICE_X18Y120_AQ),
.I3(CLBLM_L_X16Y121_SLICE_X22Y121_AQ),
.I4(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I5(CLBLM_R_X15Y120_SLICE_X20Y120_AQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555fcf05450)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.I2(CLBLM_R_X13Y120_SLICE_X19Y120_CO6),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I5(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y120_SLICE_X19Y120_AO6),
.Q(CLBLM_R_X13Y120_SLICE_X19Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05f505f530303f3f)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_DLUT (
.I0(CLBLM_R_X15Y122_SLICE_X21Y122_AQ),
.I1(CLBLM_R_X15Y121_SLICE_X20Y121_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I4(CLBLM_R_X15Y122_SLICE_X20Y122_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfadd5088fa8850)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X15Y121_SLICE_X20Y121_AQ),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(CLBLM_R_X15Y122_SLICE_X21Y122_AQ),
.I5(CLBLM_R_X15Y122_SLICE_X20Y122_AQ),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff750075ffff00ff)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_ALUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I2(LIOB33_X0Y155_IOB_X0Y155_I),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y122_SLICE_X21Y122_AQ),
.I5(CLBLM_R_X13Y121_SLICE_X19Y121_BO6),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y121_SLICE_X18Y121_AO6),
.Q(CLBLM_R_X13Y121_SLICE_X18Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h505003f35f5f03f3)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_DLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I1(CLBLM_R_X15Y121_SLICE_X21Y121_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X15Y121_SLICE_X20Y121_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_R_X15Y120_SLICE_X21Y120_AQ),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccccccf5f0f0f0)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I1(CLBLM_R_X13Y121_SLICE_X18Y121_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fafaee445050)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X15Y121_SLICE_X21Y121_AQ),
.I2(CLBLM_L_X12Y120_SLICE_X16Y120_AQ),
.I3(CLBLM_R_X15Y121_SLICE_X20Y121_BQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_R_X15Y120_SLICE_X21Y120_AQ),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33fd31fc30)
  ) CLBLM_R_X13Y121_SLICE_X18Y121_ALUT (
.I0(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y125_SLICE_X18Y125_BO6),
.I3(CLBLM_R_X15Y121_SLICE_X20Y121_BQ),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLM_R_X13Y121_SLICE_X18Y121_CO6),
.O5(CLBLM_R_X13Y121_SLICE_X18Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X18Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y121_SLICE_X19Y121_AO6),
.Q(CLBLM_R_X13Y121_SLICE_X19Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000000000)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_DO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfddffff1f11)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.I2(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(CLBLM_R_X13Y121_SLICE_X19Y121_DO6),
.I5(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_CO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h070007770f000fff)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I2(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_BO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffff220022)
  ) CLBLM_R_X13Y121_SLICE_X19Y121_ALUT (
.I0(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I2(1'b1),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I5(CLBLM_R_X13Y121_SLICE_X19Y121_CO6),
.O5(CLBLM_R_X13Y121_SLICE_X19Y121_AO5),
.O6(CLBLM_R_X13Y121_SLICE_X19Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y122_SLICE_X18Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X18Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dddd8888)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111bbbb05af05af)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I2(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I4(CLBLM_L_X12Y122_SLICE_X17Y122_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcc0fcc05440fcc)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I3(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff75ff000075ff)
  ) CLBLM_R_X13Y122_SLICE_X18Y122_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I2(LIOB33_X0Y151_IOB_X0Y152_I),
.I3(CLBLM_R_X13Y122_SLICE_X18Y122_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X18Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X18Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y122_SLICE_X19Y122_AO6),
.Q(CLBLM_R_X13Y122_SLICE_X19Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5030503f5f305f3f)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_DLUT (
.I0(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(CLBLM_R_X15Y122_SLICE_X20Y122_BQ),
.I5(CLBLM_R_X15Y123_SLICE_X21Y123_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_DO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3313ff5f0000cc4c)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I1(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I4(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_CO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefc302222fc30)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_BLUT (
.I0(CLBLM_R_X15Y122_SLICE_X20Y122_BQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I2(CLBLM_L_X12Y122_SLICE_X16Y122_AQ),
.I3(CLBLM_R_X15Y123_SLICE_X21Y123_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_AQ),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_BO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a0afafafafafaf)
  ) CLBLM_R_X13Y122_SLICE_X19Y122_ALUT (
.I0(CLBLM_L_X12Y123_SLICE_X17Y123_AQ),
.I1(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(CLBLM_R_X13Y124_SLICE_X19Y124_BO5),
.I5(CLBLM_R_X13Y122_SLICE_X19Y122_CO6),
.O5(CLBLM_R_X13Y122_SLICE_X19Y122_AO5),
.O6(CLBLM_R_X13Y122_SLICE_X19Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y123_SLICE_X18Y123_BO6),
.Q(CLBLM_R_X13Y123_SLICE_X18Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff03333f3f3)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(LIOB33_X0Y151_IOB_X0Y151_I),
.I3(CLBLM_R_X13Y123_SLICE_X18Y123_BQ),
.I4(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5d0c5dff550055)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.I4(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3e2f3e2f3f3f3e2)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_BLUT (
.I0(CLBLM_R_X13Y123_SLICE_X18Y123_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y123_SLICE_X18Y123_AQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_CO6),
.I4(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fff0ff404)
  ) CLBLM_R_X13Y123_SLICE_X18Y123_ALUT (
.I0(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I1(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.I5(CLBLM_R_X13Y123_SLICE_X18Y123_CO6),
.O5(CLBLM_R_X13Y123_SLICE_X18Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X18Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y123_SLICE_X19Y123_AO6),
.Q(CLBLM_R_X13Y123_SLICE_X19Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333ffaabbbb)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_DLUT (
.I0(LIOB33_X0Y151_IOB_X0Y151_I),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_AQ),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_DO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_CO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_BO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3e2f3e2f3f3f3e2)
  ) CLBLM_R_X13Y123_SLICE_X19Y123_ALUT (
.I0(CLBLM_R_X13Y123_SLICE_X19Y123_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I3(CLBLM_R_X13Y123_SLICE_X19Y123_BO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_AO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.O5(CLBLM_R_X13Y123_SLICE_X19Y123_AO5),
.O6(CLBLM_R_X13Y123_SLICE_X19Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y124_SLICE_X18Y124_AO6),
.Q(CLBLM_R_X13Y124_SLICE_X18Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y124_SLICE_X18Y124_BO6),
.Q(CLBLM_R_X13Y124_SLICE_X18Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddf5a08888f5a0)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X16Y125_SLICE_X22Y125_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bb050511bbafaf)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X16Y125_SLICE_X22Y125_AQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33fd31fc30)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_BLUT (
.I0(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_DO6),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AQ),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_R_X15Y123_SLICE_X20Y123_BO6),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002f2fff00ffff)
  ) CLBLM_R_X13Y124_SLICE_X18Y124_ALUT (
.I0(LIOB33_X0Y155_IOB_X0Y155_I),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I2(CLBLM_L_X16Y123_SLICE_X22Y123_AO5),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_CO6),
.O5(CLBLM_R_X13Y124_SLICE_X18Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X18Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y124_SLICE_X19Y124_AO6),
.Q(CLBLM_R_X13Y124_SLICE_X19Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff4ff000f444f)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_DLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I5(CLBLM_R_X13Y124_SLICE_X18Y124_BQ),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_DO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff4f04f0f4400)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(CLBLM_R_X13Y124_SLICE_X19Y124_AQ),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_CO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000100fffffffd)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_BO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ffdfc0d0c)
  ) CLBLM_R_X13Y124_SLICE_X19Y124_ALUT (
.I0(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.I1(CLBLM_R_X15Y124_SLICE_X20Y124_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_X0Y155_IOB_X0Y156_I),
.I4(CLBLM_L_X16Y125_SLICE_X22Y125_AQ),
.I5(CLBLM_R_X13Y124_SLICE_X19Y124_CO6),
.O5(CLBLM_R_X13Y124_SLICE_X19Y124_AO5),
.O6(CLBLM_R_X13Y124_SLICE_X19Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y125_SLICE_X18Y125_AO6),
.Q(CLBLM_R_X13Y125_SLICE_X18Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaeaa0c00aeaa)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I5(CLBLM_R_X13Y125_SLICE_X18Y125_AQ),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505f5f5010531f5)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X12Y126_SLICE_X17Y126_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I4(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000020)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfafffafa)
  ) CLBLM_R_X13Y125_SLICE_X18Y125_ALUT (
.I0(CLBLM_R_X13Y125_SLICE_X18Y125_DO6),
.I1(CLBLM_R_X13Y124_SLICE_X18Y124_AQ),
.I2(CLBLM_R_X15Y125_SLICE_X21Y125_CO5),
.I3(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X13Y125_SLICE_X18Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X18Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y125_SLICE_X19Y125_AO6),
.Q(CLBLM_R_X13Y125_SLICE_X19Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h503050305f305f30)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_DLUT (
.I0(CLBLM_R_X15Y124_SLICE_X20Y124_AQ),
.I1(CLBLM_R_X15Y125_SLICE_X21Y125_BQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y130_SLICE_X18Y130_BQ),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_DO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03f303f350505f5f)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_CLUT (
.I0(CLBLM_R_X15Y129_SLICE_X20Y129_AQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I4(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_CO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h01510b5ba1f1abfb)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X15Y125_SLICE_X21Y125_BQ),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BQ),
.I4(CLBLM_R_X15Y124_SLICE_X20Y124_AQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_BO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd8ddddddd8)
  ) CLBLM_R_X13Y125_SLICE_X19Y125_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I2(CLBLM_R_X13Y124_SLICE_X19Y124_BO6),
.I3(CLBLM_R_X15Y125_SLICE_X20Y125_AO6),
.I4(LIOB33_X0Y151_IOB_X0Y152_I),
.I5(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.O5(CLBLM_R_X13Y125_SLICE_X19Y125_AO5),
.O6(CLBLM_R_X13Y125_SLICE_X19Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y126_SLICE_X18Y126_BO6),
.Q(CLBLM_R_X13Y126_SLICE_X18Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff03333f3f3)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I2(LIOB33_X0Y151_IOB_X0Y151_I),
.I3(CLBLM_R_X13Y126_SLICE_X18Y126_BQ),
.I4(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccddccf0f0f5f0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_CLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I1(CLBLM_R_X13Y126_SLICE_X18Y126_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0f0ffee)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_BLUT (
.I0(CLBLM_R_X13Y126_SLICE_X18Y126_DO6),
.I1(CLBLM_L_X12Y126_SLICE_X17Y126_CO6),
.I2(CLBLM_L_X12Y124_SLICE_X17Y124_AQ),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3d1f3c0)
  ) CLBLM_R_X13Y126_SLICE_X18Y126_ALUT (
.I0(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y125_SLICE_X21Y125_BQ),
.I3(CLBLM_R_X13Y125_SLICE_X18Y125_BO5),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(CLBLM_R_X13Y126_SLICE_X18Y126_CO6),
.O5(CLBLM_R_X13Y126_SLICE_X18Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X18Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_AO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y126_SLICE_X19Y126_BO6),
.Q(CLBLM_R_X13Y126_SLICE_X19Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff8080ff8080)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I3(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I5(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_DO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0503553355335533)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_CLUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_BQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_CO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1f3d1f3f3f3f3)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_BLUT (
.I0(CLBLM_L_X16Y125_SLICE_X22Y125_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y126_SLICE_X19Y126_AQ),
.I3(LIOB33_X0Y155_IOB_X0Y155_I),
.I4(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I5(CLBLM_R_X13Y126_SLICE_X19Y126_CO6),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_BO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcacacfca)
  ) CLBLM_R_X13Y126_SLICE_X19Y126_ALUT (
.I0(CLBLM_R_X13Y126_SLICE_X19Y126_DO6),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(LIOB33_X0Y153_IOB_X0Y154_I),
.I4(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.I5(CLBLM_R_X15Y122_SLICE_X20Y122_CO6),
.O5(CLBLM_R_X13Y126_SLICE_X19Y126_AO5),
.O6(CLBLM_R_X13Y126_SLICE_X19Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.Q(CLBLM_R_X13Y127_SLICE_X18Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaeeeefffaffee)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_DO6),
.I1(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(LIOB33_X0Y157_IOB_X0Y157_I),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I5(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfff00f0c0f00)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_BO6),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I5(CLBLM_R_X13Y130_SLICE_X18Y130_BQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y127_SLICE_X19Y127_AO6),
.Q(CLBLM_R_X13Y127_SLICE_X19Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cf03df57df57)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_DLUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I3(CLBLM_R_X13Y127_SLICE_X19Y127_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafefafeaaeeffff)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_BLUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_CO6),
.I1(LIOB33_X0Y151_IOB_X0Y151_I),
.I2(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_DO6),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ffafe0a0e)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X19Y127_DO6),
.I1(LIOB33_X0Y151_IOB_X0Y152_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_CO6),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_BQ),
.I5(CLBLM_R_X13Y127_SLICE_X19Y127_CO6),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_BO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff303fffffbab)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_CLUT (
.I0(LIOB33_X0Y153_IOB_X0Y153_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I2(CLBLM_R_X15Y128_SLICE_X21Y128_CO6),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_DO6),
.I5(CLBLM_R_X15Y128_SLICE_X21Y128_BO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888dddd8d8d)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_BQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I3(1'b1),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000020000000)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h307530753075ffff)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_DLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000d0d0d00)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300f3f0bbaafbfa)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_AO6),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022322233)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.I2(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I3(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_BO5),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffceceffffff0a)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_CLUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_DO6),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033302220)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_BLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I4(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_AO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0cc00)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_CO6),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y129_SLICE_X19Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X19Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3333333)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y128_SLICE_X19Y128_DO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020000000000000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffb3f7a0f5)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_BLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff40f04fff40f04)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X13Y129_SLICE_X19Y129_BO6),
.I4(CLBLM_L_X12Y127_SLICE_X17Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y130_SLICE_X18Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X18Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y130_SLICE_X18Y130_BO6),
.Q(CLBLM_R_X13Y130_SLICE_X18Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef4fffffef4fef4)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_DLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_DO6),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_BQ),
.I4(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I5(LIOB33_X0Y155_IOB_X0Y156_I),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdf8f8fffdfff8)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_CLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.I3(LIOB33_X0Y155_IOB_X0Y155_I),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I5(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeaaf0f0eeaa)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_BLUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I2(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcac0cac0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_ALUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y130_SLICE_X18Y130_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X19Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffefafeeffeeaa)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_CLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I5(LIOB33_X0Y155_IOB_X0Y156_I),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33fa32aa22)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I3(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y131_SLICE_X18Y131_AO6),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X13Y131_SLICE_X18Y131_BO6),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeafffffbeafbea)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_DLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I2(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I5(LIOB33_X0Y153_IOB_X0Y154_I),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fffffff4f4f4)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_CLUT (
.I0(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I1(LIOB33_X0Y153_IOB_X0Y154_I),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_DO6),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffcca0cca0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I1(CLBLM_R_X15Y130_SLICE_X20Y130_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y131_SLICE_X18Y131_CO6),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33fa32aa22)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_ALUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_CO6),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa55ff1b1b1b1b)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X15Y126_SLICE_X21Y126_AQ),
.I2(CLBLM_R_X15Y126_SLICE_X20Y126_AQ),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfafcfa0c0afc0a0)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_BLUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.I1(CLBLM_R_X15Y126_SLICE_X20Y126_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I5(CLBLM_R_X15Y126_SLICE_X21Y126_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffaff5fffff)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeefffffeeefeeef)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_BO6),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000200002000200)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffaff00ff32)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_CLUT (
.I0(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I1(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.I4(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000200000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00400040ffff0200)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y100_SLICE_X20Y100_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y100_SLICE_X20Y100_AO6),
.Q(CLBLM_R_X15Y100_SLICE_X20Y100_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00cfcccfcc)
  ) CLBLM_R_X15Y100_SLICE_X20Y100_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y101_SLICE_X20Y101_BO5),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_R_X15Y102_SLICE_X20Y102_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.O5(CLBLM_R_X15Y100_SLICE_X20Y100_DO5),
.O6(CLBLM_R_X15Y100_SLICE_X20Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00006fcf66cc)
  ) CLBLM_R_X15Y100_SLICE_X20Y100_CLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_CO6),
.I4(CLBLM_R_X15Y101_SLICE_X20Y101_AO5),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_R_X15Y100_SLICE_X20Y100_CO5),
.O6(CLBLM_R_X15Y100_SLICE_X20Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5aa0a0a0a0)
  ) CLBLM_R_X15Y100_SLICE_X20Y100_BLUT (
.I0(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y100_SLICE_X20Y100_BO5),
.O6(CLBLM_R_X15Y100_SLICE_X20Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5f5f5e4)
  ) CLBLM_R_X15Y100_SLICE_X20Y100_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X13Y102_SLICE_X19Y102_DO6),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_DO6),
.I4(CLBLM_R_X15Y101_SLICE_X20Y101_AO6),
.I5(CLBLM_R_X15Y100_SLICE_X20Y100_CO6),
.O5(CLBLM_R_X15Y100_SLICE_X20Y100_AO5),
.O6(CLBLM_R_X15Y100_SLICE_X20Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0880000000000000)
  ) CLBLM_R_X15Y100_SLICE_X21Y100_DLUT (
.I0(CLBLM_L_X12Y100_SLICE_X17Y100_AO6),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I2(CLBLM_R_X15Y100_SLICE_X20Y100_BO5),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I5(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.O5(CLBLM_R_X15Y100_SLICE_X21Y100_DO5),
.O6(CLBLM_R_X15Y100_SLICE_X21Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000080000000)
  ) CLBLM_R_X15Y100_SLICE_X21Y100_CLUT (
.I0(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I4(CLBLM_L_X12Y101_SLICE_X17Y101_CO6),
.I5(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.O5(CLBLM_R_X15Y100_SLICE_X21Y100_CO5),
.O6(CLBLM_R_X15Y100_SLICE_X21Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h777f88807fff8000)
  ) CLBLM_R_X15Y100_SLICE_X21Y100_BLUT (
.I0(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I2(CLBLM_L_X12Y101_SLICE_X17Y101_CO6),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I4(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I5(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.O5(CLBLM_R_X15Y100_SLICE_X21Y100_BO5),
.O6(CLBLM_R_X15Y100_SLICE_X21Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y100_SLICE_X21Y100_ALUT (
.I0(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I2(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I4(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I5(CLBLM_R_X13Y100_SLICE_X18Y100_CO6),
.O5(CLBLM_R_X15Y100_SLICE_X21Y100_AO5),
.O6(CLBLM_R_X15Y100_SLICE_X21Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055f0f500aaf0fa)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_DLUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I1(1'b1),
.I2(CLBLM_R_X15Y101_SLICE_X21Y101_BO5),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I5(CLBLM_R_X15Y101_SLICE_X20Y101_BO6),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_DO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000080000000)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_CLUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I1(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I2(CLBLM_L_X12Y101_SLICE_X17Y101_BO6),
.I3(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I4(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I5(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_CO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00077887788)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_BLUT (
.I0(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I1(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_CO6),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_BO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaaf00033cc33cc)
  ) CLBLM_R_X15Y101_SLICE_X20Y101_ALUT (
.I0(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I1(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X20Y101_AO5),
.O6(CLBLM_R_X15Y101_SLICE_X20Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000080000000)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_DLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I1(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_R_X13Y101_SLICE_X19Y101_CO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(CLBLM_R_X15Y101_SLICE_X21Y101_BO6),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_DO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800800000000000)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I1(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I4(CLBLM_R_X15Y101_SLICE_X21Y101_AO6),
.I5(CLBLM_R_X13Y101_SLICE_X19Y101_BO6),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_CO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c0003cf03cf0)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I2(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I3(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_BO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800078f078f0)
  ) CLBLM_R_X15Y101_SLICE_X21Y101_ALUT (
.I0(CLBLM_R_X13Y101_SLICE_X19Y101_DO6),
.I1(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I2(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I3(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y101_SLICE_X21Y101_AO5),
.O6(CLBLM_R_X15Y101_SLICE_X21Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y102_SLICE_X20Y102_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y102_SLICE_X20Y102_AO6),
.Q(CLBLM_R_X15Y102_SLICE_X20Y102_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffccff0000cccc)
  ) CLBLM_R_X15Y102_SLICE_X20Y102_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y101_SLICE_X21Y101_AO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(CLBLM_R_X15Y102_SLICE_X20Y102_BO6),
.O5(CLBLM_R_X15Y102_SLICE_X20Y102_DO5),
.O6(CLBLM_R_X15Y102_SLICE_X20Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1717ffffe8e80000)
  ) CLBLM_R_X15Y102_SLICE_X20Y102_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_L_X12Y103_SLICE_X17Y103_CO6),
.I2(CLBLM_R_X13Y101_SLICE_X19Y101_AO5),
.I3(1'b1),
.I4(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I5(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.O5(CLBLM_R_X15Y102_SLICE_X20Y102_CO5),
.O6(CLBLM_R_X15Y102_SLICE_X20Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af078f078f0f0f0)
  ) CLBLM_R_X15Y102_SLICE_X20Y102_BLUT (
.I0(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I1(CLBLM_R_X13Y101_SLICE_X19Y101_AO5),
.I2(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_CO6),
.O5(CLBLM_R_X15Y102_SLICE_X20Y102_BO5),
.O6(CLBLM_R_X15Y102_SLICE_X20Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3e2f3e2)
  ) CLBLM_R_X15Y102_SLICE_X20Y102_ALUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I3(CLBLM_R_X15Y103_SLICE_X20Y103_BO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y101_SLICE_X20Y101_DO6),
.O5(CLBLM_R_X15Y102_SLICE_X20Y102_AO5),
.O6(CLBLM_R_X15Y102_SLICE_X20Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a55a0000a55a)
  ) CLBLM_R_X15Y102_SLICE_X21Y102_DLUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_R_X15Y102_SLICE_X21Y102_AO5),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y102_SLICE_X21Y102_DO5),
.O6(CLBLM_R_X15Y102_SLICE_X21Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hecccccccccccccc8)
  ) CLBLM_R_X15Y102_SLICE_X21Y102_CLUT (
.I0(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I5(CLBLM_L_X12Y103_SLICE_X17Y103_BO6),
.O5(CLBLM_R_X15Y102_SLICE_X21Y102_CO5),
.O6(CLBLM_R_X15Y102_SLICE_X21Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y102_SLICE_X21Y102_BLUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I1(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I2(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I3(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I4(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I5(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.O5(CLBLM_R_X15Y102_SLICE_X21Y102_BO5),
.O6(CLBLM_R_X15Y102_SLICE_X21Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaa8a8eaaaaaa8)
  ) CLBLM_R_X15Y102_SLICE_X21Y102_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_L_X12Y103_SLICE_X17Y103_BO6),
.I2(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_R_X13Y102_SLICE_X18Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y102_SLICE_X21Y102_AO5),
.O6(CLBLM_R_X15Y102_SLICE_X21Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000800000000000)
  ) CLBLM_R_X15Y103_SLICE_X20Y103_DLUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I1(CLBLM_R_X13Y103_SLICE_X19Y103_AO5),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_L_X12Y101_SLICE_X17Y101_AO6),
.I4(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I5(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.O5(CLBLM_R_X15Y103_SLICE_X20Y103_DO5),
.O6(CLBLM_R_X15Y103_SLICE_X20Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a7878f0f0f0f0f0)
  ) CLBLM_R_X15Y103_SLICE_X20Y103_CLUT (
.I0(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I1(CLBLM_R_X13Y103_SLICE_X19Y103_AO5),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_L_X12Y101_SLICE_X17Y101_AO6),
.I4(CLBLM_R_X13Y100_SLICE_X18Y100_AQ),
.I5(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.O5(CLBLM_R_X15Y103_SLICE_X20Y103_CO5),
.O6(CLBLM_R_X15Y103_SLICE_X20Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbffbbfffaffaa)
  ) CLBLM_R_X15Y103_SLICE_X20Y103_BLUT (
.I0(CLBLM_R_X15Y102_SLICE_X21Y102_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(CLBLM_R_X15Y109_SLICE_X20Y109_AO6),
.I4(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I5(CLBLM_R_X13Y102_SLICE_X19Y102_BO6),
.O5(CLBLM_R_X15Y103_SLICE_X20Y103_BO5),
.O6(CLBLM_R_X15Y103_SLICE_X20Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000007fff8000)
  ) CLBLM_R_X15Y103_SLICE_X20Y103_ALUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I1(CLBLM_R_X13Y100_SLICE_X19Y100_AO6),
.I2(CLBLM_R_X15Y102_SLICE_X20Y102_AQ),
.I3(CLBLM_R_X15Y100_SLICE_X20Y100_AQ),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y103_SLICE_X20Y103_AO5),
.O6(CLBLM_R_X15Y103_SLICE_X20Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLM_R_X15Y103_SLICE_X21Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y103_SLICE_X20Y103_AO5),
.I2(CLBLM_R_X15Y103_SLICE_X20Y103_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y103_SLICE_X21Y103_DO5),
.O6(CLBLM_R_X15Y103_SLICE_X21Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff80fe00ff80fe00)
  ) CLBLM_R_X15Y103_SLICE_X21Y103_CLUT (
.I0(CLBLM_R_X15Y102_SLICE_X21Y102_CO6),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I4(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y103_SLICE_X21Y103_CO5),
.O6(CLBLM_R_X15Y103_SLICE_X21Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbaff30)
  ) CLBLM_R_X15Y103_SLICE_X21Y103_BLUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_R_X15Y103_SLICE_X20Y103_CO6),
.I3(CLBLM_L_X16Y110_SLICE_X23Y110_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I5(CLBLM_R_X15Y103_SLICE_X21Y103_AO5),
.O5(CLBLM_R_X15Y103_SLICE_X21Y103_BO5),
.O6(CLBLM_R_X15Y103_SLICE_X21Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3021123022111122)
  ) CLBLM_R_X15Y103_SLICE_X21Y103_ALUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I3(CLBLM_R_X15Y102_SLICE_X21Y102_CO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y103_SLICE_X21Y103_AO5),
.O6(CLBLM_R_X15Y103_SLICE_X21Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y104_SLICE_X20Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y104_SLICE_X20Y104_AO6),
.Q(CLBLM_R_X15Y104_SLICE_X20Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X15Y104_SLICE_X20Y104_DLUT (
.I0(CLBLM_L_X16Y103_SLICE_X23Y103_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X15Y101_SLICE_X20Y101_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y104_SLICE_X20Y104_DO5),
.O6(CLBLM_R_X15Y104_SLICE_X20Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X15Y104_SLICE_X20Y104_CLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I4(1'b1),
.I5(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.O5(CLBLM_R_X15Y104_SLICE_X20Y104_CO5),
.O6(CLBLM_R_X15Y104_SLICE_X20Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbbfbaafa)
  ) CLBLM_R_X15Y104_SLICE_X20Y104_BLUT (
.I0(CLBLM_R_X15Y108_SLICE_X20Y108_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_R_X13Y102_SLICE_X19Y102_BO6),
.I5(CLBLM_R_X15Y109_SLICE_X20Y109_AO6),
.O5(CLBLM_R_X15Y104_SLICE_X20Y104_BO5),
.O6(CLBLM_R_X15Y104_SLICE_X20Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5a0f5e4)
  ) CLBLM_R_X15Y104_SLICE_X20Y104_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X15Y102_SLICE_X20Y102_BO6),
.I2(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I3(CLBLM_R_X15Y104_SLICE_X20Y104_BO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I5(CLBLM_R_X15Y102_SLICE_X21Y102_DO6),
.O5(CLBLM_R_X15Y104_SLICE_X20Y104_AO5),
.O6(CLBLM_R_X15Y104_SLICE_X20Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y104_SLICE_X21Y104_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y104_SLICE_X21Y104_AO6),
.Q(CLBLM_R_X15Y104_SLICE_X21Y104_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y104_SLICE_X21Y104_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y104_SLICE_X21Y104_BO6),
.Q(CLBLM_R_X15Y104_SLICE_X21Y104_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff003300550011)
  ) CLBLM_R_X15Y104_SLICE_X21Y104_DLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I1(CLBLM_L_X16Y103_SLICE_X22Y103_CO6),
.I2(1'b1),
.I3(CLBLM_R_X15Y109_SLICE_X21Y109_BO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_R_X15Y104_SLICE_X21Y104_DO5),
.O6(CLBLM_R_X15Y104_SLICE_X21Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffcfffafffe)
  ) CLBLM_R_X15Y104_SLICE_X21Y104_CLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X15Y103_SLICE_X20Y103_CO6),
.I2(CLBLM_R_X15Y108_SLICE_X21Y108_CO6),
.I3(CLBLM_L_X16Y110_SLICE_X23Y110_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_R_X15Y104_SLICE_X21Y104_CO5),
.O6(CLBLM_R_X15Y104_SLICE_X21Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffae5504)
  ) CLBLM_R_X15Y104_SLICE_X21Y104_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X15Y100_SLICE_X21Y100_BO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I3(CLBLM_R_X15Y103_SLICE_X21Y103_AO5),
.I4(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I5(CLBLM_R_X15Y104_SLICE_X21Y104_CO6),
.O5(CLBLM_R_X15Y104_SLICE_X21Y104_BO5),
.O6(CLBLM_R_X15Y104_SLICE_X21Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fb0000f3fbf3fb)
  ) CLBLM_R_X15Y104_SLICE_X21Y104_ALUT (
.I0(CLBLM_R_X15Y103_SLICE_X21Y103_DO6),
.I1(CLBLM_L_X16Y104_SLICE_X22Y104_CO6),
.I2(CLBLM_R_X15Y103_SLICE_X21Y103_AO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I4(LIOB33_X0Y193_IOB_X0Y193_I),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y104_SLICE_X21Y104_AO5),
.O6(CLBLM_R_X15Y104_SLICE_X21Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff30ba30ba)
  ) CLBLM_R_X15Y105_SLICE_X20Y105_DLUT (
.I0(CLBLM_R_X15Y105_SLICE_X21Y105_BO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(CLBLM_L_X16Y103_SLICE_X22Y103_CO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y106_SLICE_X20Y106_DO6),
.O5(CLBLM_R_X15Y105_SLICE_X20Y105_DO5),
.O6(CLBLM_R_X15Y105_SLICE_X20Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe80000000)
  ) CLBLM_R_X15Y105_SLICE_X20Y105_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I1(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.I2(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I3(CLBLM_R_X15Y102_SLICE_X21Y102_CO6),
.I4(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X15Y105_SLICE_X20Y105_CO5),
.O6(CLBLM_R_X15Y105_SLICE_X20Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000080000000)
  ) CLBLM_R_X15Y105_SLICE_X20Y105_BLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I1(CLBLM_R_X15Y101_SLICE_X20Y101_CO6),
.I2(CLBLM_R_X15Y103_SLICE_X20Y103_AO6),
.I3(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I4(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I5(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.O5(CLBLM_R_X15Y105_SLICE_X20Y105_BO5),
.O6(CLBLM_R_X15Y105_SLICE_X20Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0700080e0f0100)
  ) CLBLM_R_X15Y105_SLICE_X20Y105_ALUT (
.I0(CLBLM_L_X16Y101_SLICE_X22Y101_AQ),
.I1(CLBLM_R_X15Y102_SLICE_X21Y102_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(CLBLM_L_X16Y102_SLICE_X22Y102_AQ),
.O5(CLBLM_R_X15Y105_SLICE_X20Y105_AO5),
.O6(CLBLM_R_X15Y105_SLICE_X20Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y105_SLICE_X21Y105_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y105_SLICE_X21Y105_AO5),
.Q(CLBLM_R_X15Y105_SLICE_X21Y105_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff00ffcfffcc)
  ) CLBLM_R_X15Y105_SLICE_X21Y105_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y104_SLICE_X23Y104_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X15Y105_SLICE_X21Y105_CO6),
.I4(CLBLM_R_X15Y105_SLICE_X21Y105_BO5),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.O5(CLBLM_R_X15Y105_SLICE_X21Y105_DO5),
.O6(CLBLM_R_X15Y105_SLICE_X21Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00770f8f0f7f0088)
  ) CLBLM_R_X15Y105_SLICE_X21Y105_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I1(CLBLM_R_X15Y102_SLICE_X21Y102_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I5(CLBLM_R_X15Y104_SLICE_X20Y104_CO6),
.O5(CLBLM_R_X15Y105_SLICE_X21Y105_CO5),
.O6(CLBLM_R_X15Y105_SLICE_X21Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffaa005af0f0f0)
  ) CLBLM_R_X15Y105_SLICE_X21Y105_BLUT (
.I0(CLBLM_L_X16Y103_SLICE_X23Y103_CO6),
.I1(1'b1),
.I2(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I3(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I4(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y105_SLICE_X21Y105_BO5),
.O6(CLBLM_R_X15Y105_SLICE_X21Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000ffee00ee)
  ) CLBLM_R_X15Y105_SLICE_X21Y105_ALUT (
.I0(CLBLM_R_X15Y105_SLICE_X21Y105_DO6),
.I1(CLBLM_L_X16Y105_SLICE_X22Y105_CO6),
.I2(CLBLM_R_X15Y102_SLICE_X21Y102_BO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y105_SLICE_X21Y105_AO5),
.O6(CLBLM_R_X15Y105_SLICE_X21Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y106_SLICE_X20Y106_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y106_SLICE_X20Y106_AO6),
.Q(CLBLM_R_X15Y106_SLICE_X20Y106_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffc0dac0f0)
  ) CLBLM_R_X15Y106_SLICE_X20Y106_DLUT (
.I0(CLBLM_R_X15Y100_SLICE_X21Y100_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_L_X16Y104_SLICE_X22Y104_BQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(CLBLM_L_X16Y109_SLICE_X23Y109_BO6),
.O5(CLBLM_R_X15Y106_SLICE_X20Y106_DO5),
.O6(CLBLM_R_X15Y106_SLICE_X20Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeefeaafa)
  ) CLBLM_R_X15Y106_SLICE_X20Y106_CLUT (
.I0(CLBLM_R_X15Y105_SLICE_X20Y105_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_R_X15Y104_SLICE_X20Y104_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_L_X16Y104_SLICE_X23Y104_AQ),
.I5(CLBLM_R_X15Y109_SLICE_X20Y109_BO6),
.O5(CLBLM_R_X15Y106_SLICE_X20Y106_CO5),
.O6(CLBLM_R_X15Y106_SLICE_X20Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff22fffffff2)
  ) CLBLM_R_X15Y106_SLICE_X20Y106_BLUT (
.I0(CLBLM_R_X15Y104_SLICE_X20Y104_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I2(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I3(CLBLM_R_X15Y109_SLICE_X20Y109_BO6),
.I4(CLBLM_R_X15Y109_SLICE_X20Y109_CO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_R_X15Y106_SLICE_X20Y106_BO5),
.O6(CLBLM_R_X15Y106_SLICE_X20Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffa55515550)
  ) CLBLM_R_X15Y106_SLICE_X20Y106_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I2(CLBLM_R_X15Y105_SLICE_X20Y105_AO6),
.I3(CLBLM_R_X15Y106_SLICE_X20Y106_BO6),
.I4(CLBLM_L_X16Y105_SLICE_X23Y105_AO6),
.I5(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.O5(CLBLM_R_X15Y106_SLICE_X20Y106_AO5),
.O6(CLBLM_R_X15Y106_SLICE_X20Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3b0a3b0a)
  ) CLBLM_R_X15Y106_SLICE_X21Y106_DLUT (
.I0(CLBLM_R_X15Y106_SLICE_X21Y106_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_R_X15Y106_SLICE_X21Y106_CO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_CO5),
.O5(CLBLM_R_X15Y106_SLICE_X21Y106_DO5),
.O6(CLBLM_R_X15Y106_SLICE_X21Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h57ff7fffa8008000)
  ) CLBLM_R_X15Y106_SLICE_X21Y106_CLUT (
.I0(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I1(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I2(CLBLM_R_X15Y101_SLICE_X21Y101_DO6),
.I3(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I4(CLBLM_R_X15Y105_SLICE_X21Y105_AO6),
.I5(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.O5(CLBLM_R_X15Y106_SLICE_X21Y106_CO5),
.O6(CLBLM_R_X15Y106_SLICE_X21Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1fe0ff007f80ff00)
  ) CLBLM_R_X15Y106_SLICE_X21Y106_BLUT (
.I0(CLBLM_R_X15Y101_SLICE_X21Y101_CO6),
.I1(CLBLM_L_X16Y105_SLICE_X23Y105_AO5),
.I2(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I3(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I4(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I5(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.O5(CLBLM_R_X15Y106_SLICE_X21Y106_BO5),
.O6(CLBLM_R_X15Y106_SLICE_X21Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf708ff00ff00ef10)
  ) CLBLM_R_X15Y106_SLICE_X21Y106_ALUT (
.I0(CLBLM_R_X15Y105_SLICE_X20Y105_CO6),
.I1(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I4(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I5(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.O5(CLBLM_R_X15Y106_SLICE_X21Y106_AO5),
.O6(CLBLM_R_X15Y106_SLICE_X21Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y107_SLICE_X20Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y107_SLICE_X20Y107_AO6),
.Q(CLBLM_R_X15Y107_SLICE_X20Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heecceeccaa00aa00)
  ) CLBLM_R_X15Y107_SLICE_X20Y107_DLUT (
.I0(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I1(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X15Y107_SLICE_X20Y107_DO5),
.O6(CLBLM_R_X15Y107_SLICE_X20Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c03030c0a09060a)
  ) CLBLM_R_X15Y107_SLICE_X20Y107_CLUT (
.I0(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I1(CLBLM_R_X15Y107_SLICE_X21Y107_AO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y107_SLICE_X20Y107_CO5),
.O6(CLBLM_R_X15Y107_SLICE_X20Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc03030c0c)
  ) CLBLM_R_X15Y107_SLICE_X20Y107_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y105_SLICE_X20Y105_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I3(1'b1),
.I4(CLBLM_L_X16Y106_SLICE_X22Y106_BO5),
.I5(1'b1),
.O5(CLBLM_R_X15Y107_SLICE_X20Y107_BO5),
.O6(CLBLM_R_X15Y107_SLICE_X20Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33ff33fe32)
  ) CLBLM_R_X15Y107_SLICE_X20Y107_ALUT (
.I0(CLBLM_R_X15Y107_SLICE_X20Y107_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y107_SLICE_X20Y107_DO6),
.I3(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I4(CLBLM_L_X16Y107_SLICE_X23Y107_AO6),
.I5(CLBLM_R_X15Y107_SLICE_X20Y107_CO6),
.O5(CLBLM_R_X15Y107_SLICE_X20Y107_AO5),
.O6(CLBLM_R_X15Y107_SLICE_X20Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y107_SLICE_X21Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y107_SLICE_X21Y107_BO6),
.Q(CLBLM_R_X15Y107_SLICE_X21Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y107_SLICE_X21Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y107_SLICE_X21Y107_CO6),
.Q(CLBLM_R_X15Y107_SLICE_X21Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h22111122f2f1f1f2)
  ) CLBLM_R_X15Y107_SLICE_X21Y107_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(CLBLM_L_X16Y107_SLICE_X23Y107_DO6),
.I3(CLBLM_R_X15Y107_SLICE_X20Y107_AQ),
.I4(CLBLM_R_X15Y107_SLICE_X21Y107_AO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.O5(CLBLM_R_X15Y107_SLICE_X21Y107_DO5),
.O6(CLBLM_R_X15Y107_SLICE_X21Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaccaaffaafc)
  ) CLBLM_R_X15Y107_SLICE_X21Y107_CLUT (
.I0(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.I1(CLBLM_R_X15Y107_SLICE_X20Y107_CO5),
.I2(CLBLM_R_X15Y106_SLICE_X21Y106_BO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y108_SLICE_X21Y108_BO6),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.O5(CLBLM_R_X15Y107_SLICE_X21Y107_CO5),
.O6(CLBLM_R_X15Y107_SLICE_X21Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffaeffae)
  ) CLBLM_R_X15Y107_SLICE_X21Y107_BLUT (
.I0(CLBLM_R_X15Y107_SLICE_X21Y107_DO6),
.I1(CLBLM_R_X15Y107_SLICE_X20Y107_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_R_X15Y108_SLICE_X21Y108_DO6),
.I4(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y107_SLICE_X21Y107_BO5),
.O6(CLBLM_R_X15Y107_SLICE_X21Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ee00ffaaaa00)
  ) CLBLM_R_X15Y107_SLICE_X21Y107_ALUT (
.I0(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.I1(CLBLM_L_X16Y108_SLICE_X22Y108_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I4(CLBLM_R_X15Y105_SLICE_X20Y105_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y107_SLICE_X21Y107_AO5),
.O6(CLBLM_R_X15Y107_SLICE_X21Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h60606060ff60ff60)
  ) CLBLM_R_X15Y108_SLICE_X20Y108_DLUT (
.I0(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X15Y108_SLICE_X20Y108_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X15Y108_SLICE_X20Y108_DO5),
.O6(CLBLM_R_X15Y108_SLICE_X20Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLM_R_X15Y108_SLICE_X20Y108_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.O5(CLBLM_R_X15Y108_SLICE_X20Y108_CO5),
.O6(CLBLM_R_X15Y108_SLICE_X20Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaabaaaa)
  ) CLBLM_R_X15Y108_SLICE_X20Y108_BLUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X15Y108_SLICE_X20Y108_BO5),
.O6(CLBLM_R_X15Y108_SLICE_X20Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000000078787878)
  ) CLBLM_R_X15Y108_SLICE_X20Y108_ALUT (
.I0(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I1(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I2(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I3(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y108_SLICE_X20Y108_AO5),
.O6(CLBLM_R_X15Y108_SLICE_X20Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff555fffff000)
  ) CLBLM_R_X15Y108_SLICE_X21Y108_DLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I1(1'b1),
.I2(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I3(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I4(CLBLM_R_X15Y109_SLICE_X21Y109_DO6),
.I5(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.O5(CLBLM_R_X15Y108_SLICE_X21Y108_DO5),
.O6(CLBLM_R_X15Y108_SLICE_X21Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa0000deeecccc)
  ) CLBLM_R_X15Y108_SLICE_X21Y108_CLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X15Y110_SLICE_X21Y110_BO6),
.I2(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X15Y108_SLICE_X21Y108_CO5),
.O6(CLBLM_R_X15Y108_SLICE_X21Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff0cffae)
  ) CLBLM_R_X15Y108_SLICE_X21Y108_BLUT (
.I0(CLBLM_R_X15Y107_SLICE_X21Y107_CQ),
.I1(CLBLM_R_X15Y106_SLICE_X21Y106_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I5(CLBLM_R_X15Y109_SLICE_X21Y109_CO6),
.O5(CLBLM_R_X15Y108_SLICE_X21Y108_BO5),
.O6(CLBLM_R_X15Y108_SLICE_X21Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaabaaaa)
  ) CLBLM_R_X15Y108_SLICE_X21Y108_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X15Y108_SLICE_X21Y108_AO5),
.O6(CLBLM_R_X15Y108_SLICE_X21Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_DO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22882288ffff2288)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X15Y109_SLICE_X21Y109_AO5),
.I2(1'b1),
.I3(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I4(CLBLM_L_X16Y109_SLICE_X22Y109_CO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_CO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020002)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_BLUT (
.I0(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_BO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000030)
  ) CLBLM_R_X15Y109_SLICE_X20Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X15Y109_SLICE_X20Y109_AO5),
.O6(CLBLM_R_X15Y109_SLICE_X20Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h48484848ff48ff48)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_DLUT (
.I0(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X16Y109_SLICE_X22Y109_AO6),
.I3(CLBLM_L_X16Y109_SLICE_X23Y109_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_DO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6c0000ff6cff00)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_CLUT (
.I0(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.I1(CLBLM_R_X15Y107_SLICE_X21Y107_CQ),
.I2(CLBLM_L_X16Y109_SLICE_X22Y109_AO6),
.I3(CLBLM_L_X16Y109_SLICE_X22Y109_DO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_CO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff44f4f444)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I1(CLBLM_L_X16Y109_SLICE_X23Y109_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I4(CLBLM_R_X15Y109_SLICE_X21Y109_AO6),
.I5(CLBLM_L_X16Y109_SLICE_X23Y109_BO6),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_BO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X15Y109_SLICE_X21Y109_ALUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I2(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I3(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y109_SLICE_X21Y109_AO5),
.O6(CLBLM_R_X15Y109_SLICE_X21Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfffcccccffcc)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(CLBLM_L_X16Y109_SLICE_X23Y109_AO5),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(CLBLM_R_X15Y107_SLICE_X21Y107_BQ),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_DO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hececffecececffec)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_CLUT (
.I0(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I3(CLBLM_R_X15Y108_SLICE_X20Y108_AO5),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_CO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8100050005000500)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_BLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I2(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_CO6),
.I4(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I5(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_BO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050dc7333003300)
  ) CLBLM_R_X15Y110_SLICE_X20Y110_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I1(CLBLM_R_X15Y110_SLICE_X21Y110_BO6),
.I2(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I3(CLBLM_R_X13Y109_SLICE_X18Y109_CO6),
.I4(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X20Y110_AO5),
.O6(CLBLM_R_X15Y110_SLICE_X20Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000100)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_DLUT (
.I0(CLBLM_R_X15Y110_SLICE_X21Y110_AO6),
.I1(CLBLM_L_X16Y107_SLICE_X22Y107_AQ),
.I2(CLBLM_R_X15Y106_SLICE_X20Y106_AQ),
.I3(CLBLM_R_X15Y110_SLICE_X20Y110_BO6),
.I4(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I5(CLBLM_L_X16Y105_SLICE_X22Y105_AQ),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_DO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2211f2f155005500)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_CLUT (
.I0(CLBLM_L_X16Y109_SLICE_X22Y109_CO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I3(CLBLM_R_X15Y110_SLICE_X20Y110_BO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_CO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaa6aaa80008000)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_BLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I2(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I3(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_BO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000006ccccccc)
  ) CLBLM_R_X15Y110_SLICE_X21Y110_ALUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X15Y104_SLICE_X21Y104_AQ),
.I2(CLBLM_R_X13Y104_SLICE_X19Y104_AQ),
.I3(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I4(CLBLM_R_X15Y104_SLICE_X20Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y110_SLICE_X21Y110_AO5),
.O6(CLBLM_R_X15Y110_SLICE_X21Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2233332200000000)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I1(CLBLM_R_X15Y110_SLICE_X21Y110_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I4(CLBLM_R_X13Y115_SLICE_X18Y115_CO6),
.I5(CLBLM_R_X13Y111_SLICE_X19Y111_BO6),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_DO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0f0f0f7ffffff)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_CLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I5(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_CO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d0d050800000000)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_BLUT (
.I0(CLBLM_L_X12Y116_SLICE_X17Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_DO6),
.I3(CLBLM_R_X13Y114_SLICE_X18Y114_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I5(CLBLM_R_X15Y111_SLICE_X20Y111_CO6),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_BO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000565500003c0f)
  ) CLBLM_R_X15Y111_SLICE_X20Y111_ALUT (
.I0(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.I1(CLBLM_L_X12Y116_SLICE_X17Y116_A5Q),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_CO6),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y111_SLICE_X20Y111_AO5),
.O6(CLBLM_R_X15Y111_SLICE_X20Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y111_SLICE_X21Y111_AO6),
.Q(CLBLM_R_X15Y111_SLICE_X21Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b0a3b0a0a3b0a3b)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_DLUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I3(CLBLM_R_X15Y110_SLICE_X20Y110_AO5),
.I4(1'b1),
.I5(CLBLM_R_X15Y110_SLICE_X21Y110_AO5),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_DO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff8888ff88)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_CLUT (
.I0(CLBLM_L_X16Y104_SLICE_X22Y104_AQ),
.I1(CLBLM_L_X16Y110_SLICE_X23Y110_AO5),
.I2(1'b1),
.I3(CLBLM_L_X16Y109_SLICE_X23Y109_CO6),
.I4(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_CO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f3f5f0f5f0f7f3)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_BLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.I1(CLBLM_R_X13Y112_SLICE_X19Y112_AO6),
.I2(CLBLM_R_X15Y111_SLICE_X20Y111_AO5),
.I3(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I4(CLBLM_R_X15Y110_SLICE_X21Y110_CO5),
.I5(CLBLM_L_X16Y109_SLICE_X23Y109_CO6),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_BO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f351f351)
  ) CLBLM_R_X15Y111_SLICE_X21Y111_ALUT (
.I0(CLBLM_R_X15Y112_SLICE_X20Y112_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y197_IOB_X0Y197_I),
.I3(CLBLM_R_X15Y111_SLICE_X21Y111_BO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y111_SLICE_X21Y111_CO6),
.O5(CLBLM_R_X15Y111_SLICE_X21Y111_AO5),
.O6(CLBLM_R_X15Y111_SLICE_X21Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc54fc54f351f351)
  ) CLBLM_R_X15Y112_SLICE_X20Y112_DLUT (
.I0(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I1(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y113_SLICE_X20Y113_AO6),
.O5(CLBLM_R_X15Y112_SLICE_X20Y112_DO5),
.O6(CLBLM_R_X15Y112_SLICE_X20Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf900f9f9f900f9f9)
  ) CLBLM_R_X15Y112_SLICE_X20Y112_CLUT (
.I0(CLBLM_R_X15Y112_SLICE_X20Y112_AO6),
.I1(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y112_SLICE_X20Y112_CO5),
.O6(CLBLM_R_X15Y112_SLICE_X20Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hebbb0000ebbbebbb)
  ) CLBLM_R_X15Y112_SLICE_X20Y112_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I1(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I3(CLBLM_R_X15Y113_SLICE_X20Y113_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I5(CLBLM_L_X12Y115_SLICE_X17Y115_A5Q),
.O5(CLBLM_R_X15Y112_SLICE_X20Y112_BO5),
.O6(CLBLM_R_X15Y112_SLICE_X20Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c000c0000000)
  ) CLBLM_R_X15Y112_SLICE_X20Y112_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I2(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I3(CLBLM_R_X15Y113_SLICE_X20Y113_AO6),
.I4(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y112_SLICE_X20Y112_AO5),
.O6(CLBLM_R_X15Y112_SLICE_X20Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y112_SLICE_X21Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y112_SLICE_X21Y112_AO6),
.Q(CLBLM_R_X15Y112_SLICE_X21Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000202)
  ) CLBLM_R_X15Y112_SLICE_X21Y112_DLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.O5(CLBLM_R_X15Y112_SLICE_X21Y112_DO5),
.O6(CLBLM_R_X15Y112_SLICE_X21Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ececa0a0)
  ) CLBLM_R_X15Y112_SLICE_X21Y112_CLUT (
.I0(CLBLM_L_X16Y106_SLICE_X22Y106_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.I5(1'b1),
.O5(CLBLM_R_X15Y112_SLICE_X21Y112_CO5),
.O6(CLBLM_R_X15Y112_SLICE_X21Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020000000000003)
  ) CLBLM_R_X15Y112_SLICE_X21Y112_BLUT (
.I0(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y112_SLICE_X21Y112_BO5),
.O6(CLBLM_R_X15Y112_SLICE_X21Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffae5504ffff5555)
  ) CLBLM_R_X15Y112_SLICE_X21Y112_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X15Y110_SLICE_X21Y110_BO6),
.I2(CLBLM_R_X13Y111_SLICE_X19Y111_AO6),
.I3(CLBLM_R_X15Y112_SLICE_X21Y112_BO6),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I5(CLBLM_R_X13Y113_SLICE_X19Y113_CO6),
.O5(CLBLM_R_X15Y112_SLICE_X21Y112_AO5),
.O6(CLBLM_R_X15Y112_SLICE_X21Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_DO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_CO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_BO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X20Y113_ALUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I3(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_CO6),
.O5(CLBLM_R_X15Y113_SLICE_X20Y113_AO5),
.O6(CLBLM_R_X15Y113_SLICE_X20Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_DO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_CO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I5(CLBLM_R_X15Y114_SLICE_X21Y114_CO6),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_BO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y113_SLICE_X21Y113_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I3(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I5(CLBLM_R_X15Y115_SLICE_X21Y115_BO6),
.O5(CLBLM_R_X15Y113_SLICE_X21Y113_AO5),
.O6(CLBLM_R_X15Y113_SLICE_X21Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y114_SLICE_X20Y114_AO6),
.Q(CLBLM_R_X15Y114_SLICE_X20Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800800000000000)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_DLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_DO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888dcccc88d8cccc)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X15Y114_SLICE_X20Y114_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_R_X15Y113_SLICE_X21Y113_BO6),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_CO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_BLUT (
.I0(CLBLM_R_X15Y114_SLICE_X20Y114_DO6),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ff101f404)
  ) CLBLM_R_X15Y114_SLICE_X20Y114_ALUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I1(CLBLM_R_X15Y114_SLICE_X21Y114_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_L_X16Y114_SLICE_X23Y114_AQ),
.I4(CLBLM_L_X12Y111_SLICE_X17Y111_AQ),
.I5(CLBLM_R_X15Y114_SLICE_X20Y114_CO6),
.O5(CLBLM_R_X15Y114_SLICE_X20Y114_AO5),
.O6(CLBLM_R_X15Y114_SLICE_X20Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y114_SLICE_X21Y114_AO6),
.Q(CLBLM_R_X15Y114_SLICE_X21Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafbfafef00100040)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_L_X16Y113_SLICE_X22Y113_BO5),
.I5(CLBLM_R_X15Y114_SLICE_X21Y114_AQ),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_DO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I2(CLBLM_R_X15Y114_SLICE_X20Y114_DO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_CO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_BLUT (
.I0(CLBLM_R_X15Y115_SLICE_X21Y115_BO6),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BQ),
.I4(CLBLM_L_X12Y110_SLICE_X16Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_BO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ababff00baba)
  ) CLBLM_R_X15Y114_SLICE_X21Y114_ALUT (
.I0(CLBLM_R_X15Y114_SLICE_X21Y114_DO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X15Y112_SLICE_X21Y112_CO6),
.O5(CLBLM_R_X15Y114_SLICE_X21Y114_AO5),
.O6(CLBLM_R_X15Y114_SLICE_X21Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y115_SLICE_X20Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y115_SLICE_X20Y115_AO6),
.Q(CLBLM_R_X15Y115_SLICE_X20Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0c5ccccc0cac)
  ) CLBLM_R_X15Y115_SLICE_X20Y115_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I1(CLBLM_R_X15Y116_SLICE_X20Y116_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X15Y114_SLICE_X20Y114_BO5),
.O5(CLBLM_R_X15Y115_SLICE_X20Y115_DO5),
.O6(CLBLM_R_X15Y115_SLICE_X20Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0c0ccccc5cac)
  ) CLBLM_R_X15Y115_SLICE_X20Y115_CLUT (
.I0(CLBLM_R_X15Y114_SLICE_X20Y114_BO6),
.I1(CLBLM_R_X15Y115_SLICE_X20Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_R_X15Y115_SLICE_X20Y115_CO5),
.O6(CLBLM_R_X15Y115_SLICE_X20Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X15Y115_SLICE_X20Y115_BLUT (
.I0(CLBLM_R_X13Y113_SLICE_X19Y113_BO6),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y115_SLICE_X20Y115_BO5),
.O6(CLBLM_R_X15Y115_SLICE_X20Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33cd01ce02)
  ) CLBLM_R_X15Y115_SLICE_X20Y115_ALUT (
.I0(CLBLM_R_X15Y115_SLICE_X20Y115_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I3(CLBLM_R_X15Y116_SLICE_X20Y116_BQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I5(CLBLM_R_X15Y115_SLICE_X20Y115_CO6),
.O5(CLBLM_R_X15Y115_SLICE_X20Y115_AO5),
.O6(CLBLM_R_X15Y115_SLICE_X20Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y115_SLICE_X21Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y115_SLICE_X21Y115_AO6),
.Q(CLBLM_R_X15Y115_SLICE_X21Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y115_SLICE_X21Y115_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I5(CLBLM_R_X15Y113_SLICE_X21Y113_BO6),
.O5(CLBLM_R_X15Y115_SLICE_X21Y115_DO5),
.O6(CLBLM_R_X15Y115_SLICE_X21Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4c4c4cec4cec4c4)
  ) CLBLM_R_X15Y115_SLICE_X21Y115_CLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(CLBLM_R_X15Y115_SLICE_X21Y115_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_R_X15Y114_SLICE_X21Y114_CO6),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.O5(CLBLM_R_X15Y115_SLICE_X21Y115_CO5),
.O6(CLBLM_R_X15Y115_SLICE_X21Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y115_SLICE_X21Y115_BLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_BO6),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.O5(CLBLM_R_X15Y115_SLICE_X21Y115_BO5),
.O6(CLBLM_R_X15Y115_SLICE_X21Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a3afafa0ac)
  ) CLBLM_R_X15Y115_SLICE_X21Y115_ALUT (
.I0(CLBLM_R_X15Y115_SLICE_X20Y115_AQ),
.I1(CLBLM_R_X15Y115_SLICE_X20Y115_BO6),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I4(CLBLM_R_X15Y115_SLICE_X21Y115_CO6),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.O5(CLBLM_R_X15Y115_SLICE_X21Y115_AO5),
.O6(CLBLM_R_X15Y115_SLICE_X21Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y116_SLICE_X20Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y116_SLICE_X20Y116_AO6),
.Q(CLBLM_R_X15Y116_SLICE_X20Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y116_SLICE_X20Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y116_SLICE_X20Y116_BO6),
.Q(CLBLM_R_X15Y116_SLICE_X20Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f2ffff01020000)
  ) CLBLM_R_X15Y116_SLICE_X20Y116_DLUT (
.I0(CLBLM_R_X15Y116_SLICE_X20Y116_CO5),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(CLBLM_R_X15Y116_SLICE_X20Y116_AQ),
.O5(CLBLM_R_X15Y116_SLICE_X20Y116_DO5),
.O6(CLBLM_R_X15Y116_SLICE_X20Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800a000a000)
  ) CLBLM_R_X15Y116_SLICE_X20Y116_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X19Y113_BO6),
.I2(CLBLM_R_X15Y114_SLICE_X20Y114_DO6),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y116_SLICE_X20Y116_CO5),
.O6(CLBLM_R_X15Y116_SLICE_X20Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3d1f3d1f3c0)
  ) CLBLM_R_X15Y116_SLICE_X20Y116_BLUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y116_SLICE_X20Y116_AQ),
.I3(CLBLM_R_X15Y115_SLICE_X20Y115_DO6),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(CLBLM_R_X15Y116_SLICE_X20Y116_CO6),
.O5(CLBLM_R_X15Y116_SLICE_X20Y116_BO5),
.O6(CLBLM_R_X15Y116_SLICE_X20Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2f3e2e2f3e2)
  ) CLBLM_R_X15Y116_SLICE_X20Y116_ALUT (
.I0(CLBLM_R_X15Y116_SLICE_X20Y116_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X16Y116_SLICE_X23Y116_BQ),
.I3(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_R_X13Y113_SLICE_X19Y113_AO5),
.O5(CLBLM_R_X15Y116_SLICE_X20Y116_AO5),
.O6(CLBLM_R_X15Y116_SLICE_X20Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y116_SLICE_X21Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y116_SLICE_X21Y116_AO6),
.Q(CLBLM_R_X15Y116_SLICE_X21Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y116_SLICE_X21Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y116_SLICE_X21Y116_BO6),
.Q(CLBLM_R_X15Y116_SLICE_X21Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0a0aaaaa3aca)
  ) CLBLM_R_X15Y116_SLICE_X21Y116_DLUT (
.I0(CLBLM_R_X15Y116_SLICE_X21Y116_BQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_L_X16Y116_SLICE_X22Y116_BO5),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_R_X15Y116_SLICE_X21Y116_DO5),
.O6(CLBLM_R_X15Y116_SLICE_X21Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f44f444ff444444)
  ) CLBLM_R_X15Y116_SLICE_X21Y116_CLUT (
.I0(CLBLM_L_X16Y116_SLICE_X23Y116_DO6),
.I1(CLBLM_R_X15Y116_SLICE_X21Y116_AQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I5(CLBLM_R_X15Y113_SLICE_X21Y113_BO6),
.O5(CLBLM_R_X15Y116_SLICE_X21Y116_CO5),
.O6(CLBLM_R_X15Y116_SLICE_X21Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ef23ee22fe32)
  ) CLBLM_R_X15Y116_SLICE_X21Y116_BLUT (
.I0(CLBLM_R_X15Y116_SLICE_X21Y116_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y114_SLICE_X19Y114_AQ),
.I3(CLBLM_R_X15Y116_SLICE_X21Y116_AQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_AO5),
.O5(CLBLM_R_X15Y116_SLICE_X21Y116_BO5),
.O6(CLBLM_R_X15Y116_SLICE_X21Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333cdce0102)
  ) CLBLM_R_X15Y116_SLICE_X21Y116_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I3(CLBLM_R_X15Y113_SLICE_X21Y113_AO6),
.I4(CLBLM_R_X15Y114_SLICE_X20Y114_AQ),
.I5(CLBLM_R_X15Y116_SLICE_X21Y116_CO6),
.O5(CLBLM_R_X15Y116_SLICE_X21Y116_AO5),
.O6(CLBLM_R_X15Y116_SLICE_X21Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y117_SLICE_X20Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y117_SLICE_X20Y117_AO6),
.Q(CLBLM_R_X15Y117_SLICE_X20Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc05cccccc0acc)
  ) CLBLM_R_X15Y117_SLICE_X20Y117_DLUT (
.I0(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I1(CLBLM_R_X15Y117_SLICE_X20Y117_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X15Y117_SLICE_X20Y117_BO6),
.O5(CLBLM_R_X15Y117_SLICE_X20Y117_DO5),
.O6(CLBLM_R_X15Y117_SLICE_X20Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88aa8baa8baa88aa)
  ) CLBLM_R_X15Y117_SLICE_X20Y117_CLUT (
.I0(CLBLM_R_X15Y117_SLICE_X21Y117_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_R_X15Y117_SLICE_X20Y117_BO5),
.I5(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.O5(CLBLM_R_X15Y117_SLICE_X20Y117_CO5),
.O6(CLBLM_R_X15Y117_SLICE_X20Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X15Y117_SLICE_X20Y117_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I2(CLBLM_R_X15Y115_SLICE_X21Y115_DO6),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I4(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y117_SLICE_X20Y117_BO5),
.O6(CLBLM_R_X15Y117_SLICE_X20Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aabeaabe)
  ) CLBLM_R_X15Y117_SLICE_X20Y117_ALUT (
.I0(CLBLM_R_X15Y117_SLICE_X20Y117_DO6),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I2(CLBLM_R_X15Y118_SLICE_X20Y118_BO5),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I4(CLBLM_R_X15Y117_SLICE_X21Y117_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y117_SLICE_X20Y117_AO5),
.O6(CLBLM_R_X15Y117_SLICE_X20Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y117_SLICE_X21Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y117_SLICE_X21Y117_AO6),
.Q(CLBLM_R_X15Y117_SLICE_X21Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y117_SLICE_X21Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y117_SLICE_X21Y117_BO6),
.Q(CLBLM_R_X15Y117_SLICE_X21Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f606ff00ff00)
  ) CLBLM_R_X15Y117_SLICE_X21Y117_DLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I1(CLBLM_R_X15Y115_SLICE_X21Y115_DO6),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X15Y117_SLICE_X21Y117_BQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_R_X15Y117_SLICE_X21Y117_DO5),
.O6(CLBLM_R_X15Y117_SLICE_X21Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y117_SLICE_X21Y117_CLUT (
.I0(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I3(CLBLM_L_X16Y115_SLICE_X22Y115_BO6),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I5(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.O5(CLBLM_R_X15Y117_SLICE_X21Y117_CO5),
.O6(CLBLM_R_X15Y117_SLICE_X21Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffab00abffba00ba)
  ) CLBLM_R_X15Y117_SLICE_X21Y117_BLUT (
.I0(CLBLM_R_X15Y117_SLICE_X21Y117_DO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I2(CLBLM_L_X16Y116_SLICE_X22Y116_AO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X16Y117_SLICE_X22Y117_BQ),
.I5(CLBLM_L_X12Y111_SLICE_X17Y111_BQ),
.O5(CLBLM_R_X15Y117_SLICE_X21Y117_BO5),
.O6(CLBLM_R_X15Y117_SLICE_X21Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030fdfe3132)
  ) CLBLM_R_X15Y117_SLICE_X21Y117_ALUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y117_SLICE_X20Y117_CO6),
.I3(CLBLM_L_X16Y117_SLICE_X23Y117_AO6),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.O5(CLBLM_R_X15Y117_SLICE_X21Y117_AO5),
.O6(CLBLM_R_X15Y117_SLICE_X21Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y118_SLICE_X20Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y118_SLICE_X20Y118_AO6),
.Q(CLBLM_R_X15Y118_SLICE_X20Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y118_SLICE_X20Y118_DLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I4(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I5(CLBLM_R_X15Y115_SLICE_X21Y115_DO6),
.O5(CLBLM_R_X15Y118_SLICE_X20Y118_DO5),
.O6(CLBLM_R_X15Y118_SLICE_X20Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c8c8c8c8cdcdc8c)
  ) CLBLM_R_X15Y118_SLICE_X20Y118_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X15Y118_SLICE_X20Y118_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I4(CLBLM_R_X15Y118_SLICE_X20Y118_DO6),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_R_X15Y118_SLICE_X20Y118_CO5),
.O6(CLBLM_R_X15Y118_SLICE_X20Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_R_X15Y118_SLICE_X20Y118_BLUT (
.I0(CLBLM_R_X13Y111_SLICE_X18Y111_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I2(CLBLM_L_X16Y115_SLICE_X22Y115_BO6),
.I3(CLBLM_R_X13Y115_SLICE_X18Y115_AQ),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y118_SLICE_X20Y118_BO5),
.O6(CLBLM_R_X15Y118_SLICE_X20Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3c0c0d1e2)
  ) CLBLM_R_X15Y118_SLICE_X20Y118_ALUT (
.I0(CLBLM_R_X15Y112_SLICE_X21Y112_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y117_SLICE_X20Y117_AQ),
.I3(CLBLM_R_X15Y118_SLICE_X20Y118_BO6),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I5(CLBLM_R_X15Y118_SLICE_X20Y118_CO6),
.O5(CLBLM_R_X15Y118_SLICE_X20Y118_AO5),
.O6(CLBLM_R_X15Y118_SLICE_X20Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y118_SLICE_X21Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y118_SLICE_X21Y118_AO6),
.Q(CLBLM_R_X15Y118_SLICE_X21Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100020002000200)
  ) CLBLM_R_X15Y118_SLICE_X21Y118_DLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I5(CLBLM_L_X16Y118_SLICE_X22Y118_AO6),
.O5(CLBLM_R_X15Y118_SLICE_X21Y118_DO5),
.O6(CLBLM_R_X15Y118_SLICE_X21Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f202ff00ff00)
  ) CLBLM_R_X15Y118_SLICE_X21Y118_CLUT (
.I0(CLBLM_L_X16Y118_SLICE_X22Y118_AO6),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X15Y119_SLICE_X21Y119_BQ),
.I4(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_R_X15Y118_SLICE_X21Y118_CO5),
.O6(CLBLM_R_X15Y118_SLICE_X21Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400080008000800)
  ) CLBLM_R_X15Y118_SLICE_X21Y118_BLUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I4(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I5(CLBLM_R_X15Y119_SLICE_X21Y119_CO6),
.O5(CLBLM_R_X15Y118_SLICE_X21Y118_BO5),
.O6(CLBLM_R_X15Y118_SLICE_X21Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffe33223332)
  ) CLBLM_R_X15Y118_SLICE_X21Y118_ALUT (
.I0(CLBLM_R_X15Y118_SLICE_X21Y118_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y118_SLICE_X21Y118_AQ),
.I3(CLBLM_R_X15Y118_SLICE_X21Y118_BO6),
.I4(CLBLM_L_X16Y116_SLICE_X23Y116_DO6),
.I5(CLBLM_R_X15Y119_SLICE_X21Y119_BQ),
.O5(CLBLM_R_X15Y118_SLICE_X21Y118_AO5),
.O6(CLBLM_R_X15Y118_SLICE_X21Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y119_SLICE_X20Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y119_SLICE_X20Y119_AO6),
.Q(CLBLM_R_X15Y119_SLICE_X20Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y119_SLICE_X20Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y119_SLICE_X20Y119_DO5),
.O6(CLBLM_R_X15Y119_SLICE_X20Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc50cccccccc)
  ) CLBLM_R_X15Y119_SLICE_X20Y119_CLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I1(CLBLM_R_X15Y119_SLICE_X20Y119_AQ),
.I2(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_R_X15Y119_SLICE_X20Y119_BO5),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_R_X15Y119_SLICE_X20Y119_CO5),
.O6(CLBLM_R_X15Y119_SLICE_X20Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800aa00aa00)
  ) CLBLM_R_X15Y119_SLICE_X20Y119_BLUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I1(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y118_SLICE_X20Y118_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y119_SLICE_X20Y119_BO5),
.O6(CLBLM_R_X15Y119_SLICE_X20Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0d1f3f3c0e2)
  ) CLBLM_R_X15Y119_SLICE_X20Y119_ALUT (
.I0(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y118_SLICE_X20Y118_AQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I4(CLBLM_R_X15Y119_SLICE_X20Y119_CO6),
.I5(CLBLM_R_X15Y117_SLICE_X21Y117_CO6),
.O5(CLBLM_R_X15Y119_SLICE_X20Y119_AO5),
.O6(CLBLM_R_X15Y119_SLICE_X20Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y119_SLICE_X21Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y119_SLICE_X21Y119_AO6),
.Q(CLBLM_R_X15Y119_SLICE_X21Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y119_SLICE_X21Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y119_SLICE_X21Y119_BO6),
.Q(CLBLM_R_X15Y119_SLICE_X21Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d88d8cccccccc)
  ) CLBLM_R_X15Y119_SLICE_X21Y119_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X15Y119_SLICE_X21Y119_AQ),
.I2(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I4(CLBLM_L_X16Y119_SLICE_X22Y119_CO6),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.O5(CLBLM_R_X15Y119_SLICE_X21Y119_DO5),
.O6(CLBLM_R_X15Y119_SLICE_X21Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X15Y119_SLICE_X21Y119_CLUT (
.I0(CLBLM_R_X15Y111_SLICE_X21Y111_AQ),
.I1(CLBLM_R_X15Y117_SLICE_X21Y117_CO6),
.I2(CLBLM_L_X16Y111_SLICE_X23Y111_AQ),
.I3(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.I4(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y119_SLICE_X21Y119_CO5),
.O6(CLBLM_R_X15Y119_SLICE_X21Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0d1f3f3d1c0)
  ) CLBLM_R_X15Y119_SLICE_X21Y119_BLUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y119_SLICE_X21Y119_AQ),
.I3(CLBLM_L_X16Y111_SLICE_X22Y111_AQ),
.I4(CLBLM_R_X15Y118_SLICE_X21Y118_CO6),
.I5(CLBLM_R_X15Y119_SLICE_X21Y119_CO6),
.O5(CLBLM_R_X15Y119_SLICE_X21Y119_BO5),
.O6(CLBLM_R_X15Y119_SLICE_X21Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0bbf0bbf0aa)
  ) CLBLM_R_X15Y119_SLICE_X21Y119_ALUT (
.I0(CLBLM_R_X15Y119_SLICE_X21Y119_DO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.I2(CLBLM_L_X16Y119_SLICE_X22Y119_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y119_SLICE_X21Y119_CO5),
.I5(CLBLM_L_X16Y111_SLICE_X22Y111_BQ),
.O5(CLBLM_R_X15Y119_SLICE_X21Y119_AO5),
.O6(CLBLM_R_X15Y119_SLICE_X21Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y120_SLICE_X20Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y120_SLICE_X20Y120_AO6),
.Q(CLBLM_R_X15Y120_SLICE_X20Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y120_SLICE_X20Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y120_SLICE_X20Y120_DO5),
.O6(CLBLM_R_X15Y120_SLICE_X20Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_R_X15Y120_SLICE_X20Y120_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X15Y120_SLICE_X20Y120_CO5),
.O6(CLBLM_R_X15Y120_SLICE_X20Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0fffff8f08800)
  ) CLBLM_R_X15Y120_SLICE_X20Y120_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y120_SLICE_X20Y120_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I4(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.O5(CLBLM_R_X15Y120_SLICE_X20Y120_BO5),
.O6(CLBLM_R_X15Y120_SLICE_X20Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff40f0f0f04)
  ) CLBLM_R_X15Y120_SLICE_X20Y120_ALUT (
.I0(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I1(LIOB33_X0Y155_IOB_X0Y155_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(CLBLM_R_X15Y120_SLICE_X20Y120_BO6),
.I4(CLBLM_R_X15Y123_SLICE_X21Y123_BO6),
.I5(CLBLM_R_X15Y121_SLICE_X20Y121_AQ),
.O5(CLBLM_R_X15Y120_SLICE_X20Y120_AO5),
.O6(CLBLM_R_X15Y120_SLICE_X20Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y120_SLICE_X21Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y120_SLICE_X21Y120_AO6),
.Q(CLBLM_R_X15Y120_SLICE_X21Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y120_SLICE_X21Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y120_SLICE_X21Y120_DO5),
.O6(CLBLM_R_X15Y120_SLICE_X21Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y120_SLICE_X21Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y120_SLICE_X21Y120_CO5),
.O6(CLBLM_R_X15Y120_SLICE_X21Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080800002000)
  ) CLBLM_R_X15Y120_SLICE_X21Y120_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X15Y120_SLICE_X21Y120_BO5),
.O6(CLBLM_R_X15Y120_SLICE_X21Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0aaee)
  ) CLBLM_R_X15Y120_SLICE_X21Y120_ALUT (
.I0(CLBLM_R_X15Y120_SLICE_X21Y120_BO5),
.I1(LIOB33_X0Y155_IOB_X0Y156_I),
.I2(CLBLM_R_X13Y120_SLICE_X19Y120_AQ),
.I3(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X15Y121_SLICE_X21Y121_CO6),
.O5(CLBLM_R_X15Y120_SLICE_X21Y120_AO5),
.O6(CLBLM_R_X15Y120_SLICE_X21Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y121_SLICE_X20Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y121_SLICE_X20Y121_AO6),
.Q(CLBLM_R_X15Y121_SLICE_X20Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y121_SLICE_X20Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y121_SLICE_X20Y121_BO6),
.Q(CLBLM_R_X15Y121_SLICE_X20Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffceffffffceff0a)
  ) CLBLM_R_X15Y121_SLICE_X20Y121_DLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_R_X15Y121_SLICE_X20Y121_AQ),
.I2(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I3(CLBLM_R_X15Y120_SLICE_X20Y120_CO6),
.I4(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.O5(CLBLM_R_X15Y121_SLICE_X20Y121_DO5),
.O6(CLBLM_R_X15Y121_SLICE_X20Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000007f7f7f007f)
  ) CLBLM_R_X15Y121_SLICE_X20Y121_CLUT (
.I0(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.I5(CLBLM_R_X15Y121_SLICE_X20Y121_BQ),
.O5(CLBLM_R_X15Y121_SLICE_X20Y121_CO5),
.O6(CLBLM_R_X15Y121_SLICE_X20Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10ff33ff33ff33)
  ) CLBLM_R_X15Y121_SLICE_X20Y121_BLUT (
.I0(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_R_X15Y120_SLICE_X20Y120_AQ),
.I4(CLBLM_R_X15Y124_SLICE_X20Y124_BO5),
.I5(CLBLM_R_X15Y121_SLICE_X20Y121_CO6),
.O5(CLBLM_R_X15Y121_SLICE_X20Y121_BO5),
.O6(CLBLM_R_X15Y121_SLICE_X20Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccaaccfaccaa)
  ) CLBLM_R_X15Y121_SLICE_X20Y121_ALUT (
.I0(CLBLM_R_X15Y121_SLICE_X20Y121_DO6),
.I1(CLBLM_R_X15Y123_SLICE_X20Y123_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y121_SLICE_X20Y121_AO5),
.O6(CLBLM_R_X15Y121_SLICE_X20Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y121_SLICE_X21Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y121_SLICE_X21Y121_AO6),
.Q(CLBLM_R_X15Y121_SLICE_X21Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd555eaaac000)
  ) CLBLM_R_X15Y121_SLICE_X21Y121_DLUT (
.I0(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X15Y121_SLICE_X21Y121_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.O5(CLBLM_R_X15Y121_SLICE_X21Y121_DO5),
.O6(CLBLM_R_X15Y121_SLICE_X21Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafcccaaaacccc)
  ) CLBLM_R_X15Y121_SLICE_X21Y121_CLUT (
.I0(CLBLM_R_X15Y120_SLICE_X21Y120_AQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I4(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O5(CLBLM_R_X15Y121_SLICE_X21Y121_CO5),
.O6(CLBLM_R_X15Y121_SLICE_X21Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff88f88fff00f00)
  ) CLBLM_R_X15Y121_SLICE_X21Y121_BLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I4(CLBLM_L_X16Y121_SLICE_X22Y121_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_R_X15Y121_SLICE_X21Y121_BO5),
.O6(CLBLM_R_X15Y121_SLICE_X21Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33ee22fe32)
  ) CLBLM_R_X15Y121_SLICE_X21Y121_ALUT (
.I0(CLBLM_R_X15Y121_SLICE_X21Y121_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_L_X16Y121_SLICE_X22Y121_AQ),
.I4(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.I5(CLBLM_R_X15Y124_SLICE_X20Y124_CO6),
.O5(CLBLM_R_X15Y121_SLICE_X21Y121_AO5),
.O6(CLBLM_R_X15Y121_SLICE_X21Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y122_SLICE_X20Y122_AO6),
.Q(CLBLM_R_X15Y122_SLICE_X20Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y122_SLICE_X20Y122_BO6),
.Q(CLBLM_R_X15Y122_SLICE_X20Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h45cf55ff45005500)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_DLUT (
.I0(CLBLM_R_X15Y122_SLICE_X20Y122_BQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I3(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_DO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000020)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_CO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddff1133fdff3133)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_BLUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_BO5),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y153_IOB_X0Y153_I),
.I3(CLBLM_R_X15Y122_SLICE_X20Y122_DO6),
.I4(CLBLM_R_X13Y122_SLICE_X19Y122_AQ),
.I5(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_BO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccaaccffccfa)
  ) CLBLM_R_X15Y122_SLICE_X20Y122_ALUT (
.I0(CLBLM_R_X15Y122_SLICE_X21Y122_CO6),
.I1(CLBLM_R_X15Y122_SLICE_X20Y122_BQ),
.I2(LIOB33_X0Y153_IOB_X0Y154_I),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y122_SLICE_X20Y122_CO5),
.I5(CLBLM_L_X16Y123_SLICE_X22Y123_BO6),
.O5(CLBLM_R_X15Y122_SLICE_X20Y122_AO5),
.O6(CLBLM_R_X15Y122_SLICE_X20Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y122_SLICE_X21Y122_AO6),
.Q(CLBLM_R_X15Y122_SLICE_X21Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_DLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_DO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf8bb88bb88bb88)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_CLUT (
.I0(CLBLM_R_X15Y122_SLICE_X20Y122_AQ),
.I1(CLBLM_L_X16Y125_SLICE_X23Y125_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_CO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfafaffbbffaa)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_BLUT (
.I0(CLBLM_R_X15Y122_SLICE_X21Y122_DO6),
.I1(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.I2(CLBLM_R_X15Y122_SLICE_X21Y122_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_BO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffc0ffc0)
  ) CLBLM_R_X15Y122_SLICE_X21Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_AO6),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I3(CLBLM_R_X15Y122_SLICE_X21Y122_BO6),
.I4(CLBLM_R_X15Y123_SLICE_X21Y123_AQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y122_SLICE_X21Y122_AO5),
.O6(CLBLM_R_X15Y122_SLICE_X21Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y123_SLICE_X20Y123_AO6),
.Q(CLBLM_R_X15Y123_SLICE_X20Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0f0f0f88cccccc)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_DO6),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_DO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbffffffefffff)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_CO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00800000fffffffb)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_BO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f07755ffff)
  ) CLBLM_R_X15Y123_SLICE_X20Y123_ALUT (
.I0(CLBLM_R_X15Y123_SLICE_X20Y123_DO6),
.I1(CLBLM_L_X16Y125_SLICE_X22Y125_DO6),
.I2(CLBLM_R_X13Y121_SLICE_X19Y121_AQ),
.I3(LIOB33_X0Y153_IOB_X0Y153_I),
.I4(CLBLM_R_X15Y123_SLICE_X20Y123_CO5),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y123_SLICE_X20Y123_AO5),
.O6(CLBLM_R_X15Y123_SLICE_X20Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y123_SLICE_X21Y123_AO6),
.Q(CLBLM_R_X15Y123_SLICE_X21Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c085f0a5f0a5f0a)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_DLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_CO6),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I2(CLBLM_R_X15Y123_SLICE_X21Y123_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_DO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffdffff)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_CO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000020)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_BO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f0fff0ddf0ff)
  ) CLBLM_R_X15Y123_SLICE_X21Y123_ALUT (
.I0(CLBLM_R_X15Y123_SLICE_X21Y123_DO6),
.I1(LIOB33_X0Y153_IOB_X0Y153_I),
.I2(CLBLM_R_X13Y122_SLICE_X18Y122_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X15Y123_SLICE_X21Y123_CO5),
.I5(CLBLM_L_X12Y123_SLICE_X17Y123_CO6),
.O5(CLBLM_R_X15Y123_SLICE_X21Y123_AO5),
.O6(CLBLM_R_X15Y123_SLICE_X21Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y124_SLICE_X20Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y124_SLICE_X20Y124_AO6),
.Q(CLBLM_R_X15Y124_SLICE_X20Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeaaac000eaaa)
  ) CLBLM_R_X15Y124_SLICE_X20Y124_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I5(CLBLM_R_X15Y124_SLICE_X20Y124_AQ),
.O5(CLBLM_R_X15Y124_SLICE_X20Y124_DO5),
.O6(CLBLM_R_X15Y124_SLICE_X20Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002010000000)
  ) CLBLM_R_X15Y124_SLICE_X20Y124_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X15Y124_SLICE_X20Y124_CO5),
.O6(CLBLM_R_X15Y124_SLICE_X20Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000fbffffff)
  ) CLBLM_R_X15Y124_SLICE_X20Y124_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y124_SLICE_X20Y124_BO5),
.O6(CLBLM_R_X15Y124_SLICE_X20Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ee22ff33fe32)
  ) CLBLM_R_X15Y124_SLICE_X20Y124_ALUT (
.I0(CLBLM_R_X15Y124_SLICE_X20Y124_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_R_X15Y127_SLICE_X20Y127_AQ),
.I4(CLBLM_R_X15Y124_SLICE_X20Y124_CO5),
.I5(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.O5(CLBLM_R_X15Y124_SLICE_X20Y124_AO5),
.O6(CLBLM_R_X15Y124_SLICE_X20Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y124_SLICE_X21Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y124_SLICE_X21Y124_AO6),
.Q(CLBLM_R_X15Y124_SLICE_X21Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0faaff080c88cc)
  ) CLBLM_R_X15Y124_SLICE_X21Y124_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I3(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.O5(CLBLM_R_X15Y124_SLICE_X21Y124_DO5),
.O6(CLBLM_R_X15Y124_SLICE_X21Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff40ffff404040)
  ) CLBLM_R_X15Y124_SLICE_X21Y124_CLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.I4(CLBLM_R_X15Y125_SLICE_X21Y125_BQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.O5(CLBLM_R_X15Y124_SLICE_X21Y124_CO5),
.O6(CLBLM_R_X15Y124_SLICE_X21Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0f0e0feeff0000)
  ) CLBLM_R_X15Y124_SLICE_X21Y124_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I2(CLBLM_R_X15Y124_SLICE_X21Y124_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I5(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.O5(CLBLM_R_X15Y124_SLICE_X21Y124_BO5),
.O6(CLBLM_R_X15Y124_SLICE_X21Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1f3c0f3f3f3f3f3)
  ) CLBLM_R_X15Y124_SLICE_X21Y124_ALUT (
.I0(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I3(CLBLM_R_X15Y124_SLICE_X21Y124_BO6),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_R_X15Y123_SLICE_X21Y123_CO6),
.O5(CLBLM_R_X15Y124_SLICE_X21Y124_AO5),
.O6(CLBLM_R_X15Y124_SLICE_X21Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303f3f05050505)
  ) CLBLM_R_X15Y125_SLICE_X20Y125_DLUT (
.I0(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I1(CLBLM_R_X15Y126_SLICE_X20Y126_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(1'b1),
.I4(CLBLM_R_X15Y124_SLICE_X21Y124_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_R_X15Y125_SLICE_X20Y125_DO5),
.O6(CLBLM_R_X15Y125_SLICE_X20Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050505050303f3f3)
  ) CLBLM_R_X15Y125_SLICE_X20Y125_CLUT (
.I0(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_R_X15Y125_SLICE_X20Y125_CO5),
.O6(CLBLM_R_X15Y125_SLICE_X20Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a5f5f11bb11bb)
  ) CLBLM_R_X15Y125_SLICE_X20Y125_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I1(CLBLM_R_X15Y124_SLICE_X21Y124_AQ),
.I2(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I3(CLBLM_R_X15Y126_SLICE_X20Y126_BQ),
.I4(CLBLM_R_X15Y130_SLICE_X20Y130_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_R_X15Y125_SLICE_X20Y125_BO5),
.O6(CLBLM_R_X15Y125_SLICE_X20Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff0055aeff0c5d)
  ) CLBLM_R_X15Y125_SLICE_X20Y125_ALUT (
.I0(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I4(CLBLM_R_X13Y125_SLICE_X19Y125_AQ),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.O5(CLBLM_R_X15Y125_SLICE_X20Y125_AO5),
.O6(CLBLM_R_X15Y125_SLICE_X20Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y125_SLICE_X21Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y125_SLICE_X21Y125_AO6),
.Q(CLBLM_R_X15Y125_SLICE_X21Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y125_SLICE_X21Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y125_SLICE_X21Y125_BO6),
.Q(CLBLM_R_X15Y125_SLICE_X21Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff40ffffff404040)
  ) CLBLM_R_X15Y125_SLICE_X21Y125_DLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X15Y125_SLICE_X21Y125_AQ),
.I4(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.O5(CLBLM_R_X15Y125_SLICE_X21Y125_DO5),
.O6(CLBLM_R_X15Y125_SLICE_X21Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000008000)
  ) CLBLM_R_X15Y125_SLICE_X21Y125_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y125_SLICE_X21Y125_CO5),
.O6(CLBLM_R_X15Y125_SLICE_X21Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbbbb88bbb8)
  ) CLBLM_R_X15Y125_SLICE_X21Y125_BLUT (
.I0(CLBLM_R_X15Y125_SLICE_X21Y125_AQ),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(CLBLM_R_X15Y124_SLICE_X21Y124_CO6),
.I4(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.I5(CLBLM_R_X15Y125_SLICE_X21Y125_CO6),
.O5(CLBLM_R_X15Y125_SLICE_X21Y125_BO5),
.O6(CLBLM_R_X15Y125_SLICE_X21Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfafaccccfffa)
  ) CLBLM_R_X15Y125_SLICE_X21Y125_ALUT (
.I0(CLBLM_R_X15Y125_SLICE_X21Y125_DO6),
.I1(CLBLM_R_X15Y126_SLICE_X21Y126_AQ),
.I2(CLBLM_R_X15Y123_SLICE_X21Y123_BO5),
.I3(LIOB33_X0Y155_IOB_X0Y155_I),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.O5(CLBLM_R_X15Y125_SLICE_X21Y125_AO5),
.O6(CLBLM_R_X15Y125_SLICE_X21Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y126_SLICE_X20Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y126_SLICE_X20Y126_AO6),
.Q(CLBLM_R_X15Y126_SLICE_X20Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y126_SLICE_X20Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y126_SLICE_X20Y126_BO6),
.Q(CLBLM_R_X15Y126_SLICE_X20Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777444407770444)
  ) CLBLM_R_X15Y126_SLICE_X20Y126_DLUT (
.I0(CLBLM_R_X15Y126_SLICE_X20Y126_BQ),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O5(CLBLM_R_X15Y126_SLICE_X20Y126_DO5),
.O6(CLBLM_R_X15Y126_SLICE_X20Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff8080ff8080)
  ) CLBLM_R_X15Y126_SLICE_X20Y126_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I5(CLBLM_R_X15Y126_SLICE_X20Y126_AQ),
.O5(CLBLM_R_X15Y126_SLICE_X20Y126_CO5),
.O6(CLBLM_R_X15Y126_SLICE_X20Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffdfdf13331313)
  ) CLBLM_R_X15Y126_SLICE_X20Y126_BLUT (
.I0(CLBLM_R_X15Y126_SLICE_X20Y126_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y123_SLICE_X20Y123_CO6),
.I3(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_R_X15Y129_SLICE_X20Y129_AQ),
.O5(CLBLM_R_X15Y126_SLICE_X20Y126_BO5),
.O6(CLBLM_R_X15Y126_SLICE_X20Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffccffcc50)
  ) CLBLM_R_X15Y126_SLICE_X20Y126_ALUT (
.I0(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I1(CLBLM_R_X15Y126_SLICE_X20Y126_BQ),
.I2(LIOB33_X0Y153_IOB_X0Y154_I),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_L_X16Y126_SLICE_X22Y126_BO5),
.I5(CLBLM_R_X15Y126_SLICE_X20Y126_CO6),
.O5(CLBLM_R_X15Y126_SLICE_X20Y126_AO5),
.O6(CLBLM_R_X15Y126_SLICE_X20Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y126_SLICE_X21Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y126_SLICE_X21Y126_AO6),
.Q(CLBLM_R_X15Y126_SLICE_X21Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff02ffffff02)
  ) CLBLM_R_X15Y126_SLICE_X21Y126_DLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y126_SLICE_X21Y126_CO6),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I5(1'b1),
.O5(CLBLM_R_X15Y126_SLICE_X21Y126_DO5),
.O6(CLBLM_R_X15Y126_SLICE_X21Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ddd0ddd00000ddd)
  ) CLBLM_R_X15Y126_SLICE_X21Y126_CLUT (
.I0(CLBLM_L_X16Y126_SLICE_X23Y126_AO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X16Y126_SLICE_X23Y126_AO5),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.O5(CLBLM_R_X15Y126_SLICE_X21Y126_CO5),
.O6(CLBLM_R_X15Y126_SLICE_X21Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88fbf8bb88bb88)
  ) CLBLM_R_X15Y126_SLICE_X21Y126_BLUT (
.I0(CLBLM_R_X15Y126_SLICE_X21Y126_AQ),
.I1(CLBLM_L_X16Y125_SLICE_X23Y125_CO6),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_R_X15Y126_SLICE_X21Y126_BO5),
.O6(CLBLM_R_X15Y126_SLICE_X21Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ffdc3310)
  ) CLBLM_R_X15Y126_SLICE_X21Y126_ALUT (
.I0(CLBLM_R_X15Y126_SLICE_X21Y126_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(LIOB33_X0Y153_IOB_X0Y154_I),
.I3(CLBLM_R_X15Y126_SLICE_X21Y126_BO6),
.I4(CLBLM_R_X15Y124_SLICE_X21Y124_AQ),
.I5(CLBLM_R_X15Y129_SLICE_X21Y129_AO6),
.O5(CLBLM_R_X15Y126_SLICE_X21Y126_AO5),
.O6(CLBLM_R_X15Y126_SLICE_X21Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y127_SLICE_X20Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y127_SLICE_X20Y127_AO6),
.Q(CLBLM_R_X15Y127_SLICE_X20Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd00000ddd0ddd0)
  ) CLBLM_R_X15Y127_SLICE_X20Y127_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X16Y126_SLICE_X23Y126_BO5),
.I2(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.O5(CLBLM_R_X15Y127_SLICE_X20Y127_DO5),
.O6(CLBLM_R_X15Y127_SLICE_X20Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X15Y127_SLICE_X20Y127_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O5(CLBLM_R_X15Y127_SLICE_X20Y127_CO5),
.O6(CLBLM_R_X15Y127_SLICE_X20Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffe4ffe4e4)
  ) CLBLM_R_X15Y127_SLICE_X20Y127_BLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I2(CLBLM_R_X15Y127_SLICE_X20Y127_AQ),
.I3(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I4(LIOB33_X0Y155_IOB_X0Y155_I),
.I5(CLBLM_R_X15Y127_SLICE_X20Y127_CO6),
.O5(CLBLM_R_X15Y127_SLICE_X20Y127_BO5),
.O6(CLBLM_R_X15Y127_SLICE_X20Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f0ff00)
  ) CLBLM_R_X15Y127_SLICE_X20Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I2(CLBLM_R_X15Y126_SLICE_X20Y126_AQ),
.I3(CLBLM_R_X15Y127_SLICE_X20Y127_BO6),
.I4(LIOB33_X0Y187_IOB_X0Y187_I),
.I5(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.O5(CLBLM_R_X15Y127_SLICE_X20Y127_AO5),
.O6(CLBLM_R_X15Y127_SLICE_X20Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0003000a0002)
  ) CLBLM_R_X15Y127_SLICE_X21Y127_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I2(CLBLM_R_X15Y128_SLICE_X21Y128_AO5),
.I3(CLBLM_R_X15Y127_SLICE_X21Y127_AO5),
.I4(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I5(CLBLM_L_X16Y126_SLICE_X23Y126_BO6),
.O5(CLBLM_R_X15Y127_SLICE_X21Y127_DO5),
.O6(CLBLM_R_X15Y127_SLICE_X21Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfcfcfcfcfcfc)
  ) CLBLM_R_X15Y127_SLICE_X21Y127_CLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I2(CLBLM_R_X15Y127_SLICE_X20Y127_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_R_X15Y127_SLICE_X21Y127_CO5),
.O6(CLBLM_R_X15Y127_SLICE_X21Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff0023)
  ) CLBLM_R_X15Y127_SLICE_X21Y127_BLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I2(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I3(CLBLM_R_X15Y128_SLICE_X21Y128_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_R_X15Y127_SLICE_X21Y127_AO5),
.O5(CLBLM_R_X15Y127_SLICE_X21Y127_BO5),
.O6(CLBLM_R_X15Y127_SLICE_X21Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800200000)
  ) CLBLM_R_X15Y127_SLICE_X21Y127_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y127_SLICE_X21Y127_AO5),
.O6(CLBLM_R_X15Y127_SLICE_X21Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c0f080a)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_DLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_BO6),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_DO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf8affaaffaaffaa)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y128_SLICE_X20Y128_AO5),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_CO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000008000)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_BO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff5ff4ffffff)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_AO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7575ff753030ff30)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_DLUT (
.I0(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I1(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_DO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505000501010001)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_CLUT (
.I0(CLBLM_R_X15Y128_SLICE_X21Y128_AO6),
.I1(CLBLM_R_X15Y120_SLICE_X21Y120_BO6),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_BO5),
.I3(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I5(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_CO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5d55ffff5575)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_BLUT (
.I0(CLBLM_R_X15Y128_SLICE_X21Y128_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_BO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000004000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_AO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y129_SLICE_X20Y129_AO6),
.Q(CLBLM_R_X15Y129_SLICE_X20Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_DLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_DO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_CLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_CO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff737f505)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.I3(CLBLM_R_X15Y129_SLICE_X20Y129_AQ),
.I4(LIOB33_X0Y151_IOB_X0Y152_I),
.I5(CLBLM_R_X15Y129_SLICE_X20Y129_CO6),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_BO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ffcc)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y132_SLICE_X19Y132_AO6),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I3(CLBLM_R_X15Y129_SLICE_X20Y129_BO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_AO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeeeeeeefeeeeee)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_DLUT (
.I0(CLBLM_R_X15Y129_SLICE_X21Y129_CO6),
.I1(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_DO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefffffffeffff)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_CLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_CO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f5ffff)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X13Y114_SLICE_X19Y114_BO6),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X13Y111_SLICE_X18Y111_BO5),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_BO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000001000000)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_AO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y130_SLICE_X20Y130_AO6),
.Q(CLBLM_R_X15Y130_SLICE_X20Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y130_SLICE_X20Y130_BO6),
.Q(CLBLM_R_X15Y130_SLICE_X20Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf1fbf1fffffbf1)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_DLUT (
.I0(CLBLM_R_X13Y128_SLICE_X19Y128_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I2(CLBLM_R_X15Y130_SLICE_X21Y130_DO6),
.I3(CLBLM_R_X15Y130_SLICE_X20Y130_BQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_DO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffceffffffceff0a)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_CLUT (
.I0(LIOB33_X0Y155_IOB_X0Y155_I),
.I1(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I3(CLBLM_R_X15Y129_SLICE_X20Y129_DO6),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_CO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeee22332222)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_BLUT (
.I0(CLBLM_R_X15Y130_SLICE_X20Y130_DO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(1'b1),
.I3(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I4(LIOB33_X0Y153_IOB_X0Y153_I),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_BO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaac0aac0)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_ALUT (
.I0(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(1'b1),
.I5(CLBLM_R_X15Y130_SLICE_X20Y130_CO6),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_AO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y130_SLICE_X21Y130_AO6),
.Q(CLBLM_R_X15Y130_SLICE_X21Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_DO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff0c5d5d)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_CLUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I1(LIOB33_X0Y153_IOB_X0Y153_I),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I3(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_CO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_BO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f351f300)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_R_X15Y130_SLICE_X21Y130_BO6),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I5(CLBLM_R_X15Y130_SLICE_X21Y130_CO6),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_AO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_BO5),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_AO6),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_BO6),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000055cc000f5f)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_AQ),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_DO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000e2c0aa77)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_BQ),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_CO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00e2e2e2e2)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_BO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_CO5),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_BO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_ALUT (
.I0(LIOB33_X0Y187_IOB_X0Y187_I),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_DO5),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_AO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_AO5),
.Q(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y131_SLICE_X21Y131_AO6),
.Q(CLBLM_R_X15Y131_SLICE_X21Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.Q(CLBLM_R_X15Y131_SLICE_X21Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_DO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_CO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff0ddf088)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_CO6),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_AQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X20Y131_DO6),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_BO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfdec31313120)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_CO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_AQ),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(CLBLM_R_X15Y132_SLICE_X21Y132_DQ),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_AO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_DO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_CO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_BO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y132_SLICE_X20Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y132_SLICE_X20Y132_AO5),
.O6(CLBLM_R_X15Y132_SLICE_X20Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y132_SLICE_X21Y132_AO6),
.Q(CLBLM_R_X15Y132_SLICE_X21Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y132_SLICE_X21Y132_BO6),
.Q(CLBLM_R_X15Y132_SLICE_X21Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y132_SLICE_X21Y132_CO6),
.Q(CLBLM_R_X15Y132_SLICE_X21Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y185_IOB_X0Y186_I),
.D(CLBLM_R_X15Y132_SLICE_X21Y132_DO6),
.Q(CLBLM_R_X15Y132_SLICE_X21Y132_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfa50ff00)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X15Y132_SLICE_X21Y132_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_AQ),
.I3(CLBLM_R_X15Y132_SLICE_X21Y132_DQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_DO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00dcdc8c8c)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_R_X15Y132_SLICE_X21Y132_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I3(CLBLM_R_X15Y132_SLICE_X21Y132_BQ),
.I4(CLBLM_R_X15Y131_SLICE_X20Y131_BQ),
.I5(LIOB33_X0Y187_IOB_X0Y187_I),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_CO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffe400cc00e4)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(CLBLM_R_X15Y132_SLICE_X21Y132_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_BQ),
.I3(LIOB33_X0Y187_IOB_X0Y187_I),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(CLBLM_R_X15Y132_SLICE_X21Y132_AQ),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_BO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd3331ccec0020)
  ) CLBLM_R_X15Y132_SLICE_X21Y132_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_B5Q),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I4(CLBLM_R_X15Y118_SLICE_X21Y118_AQ),
.I5(CLBLM_R_X15Y132_SLICE_X21Y132_AQ),
.O5(CLBLM_R_X15Y132_SLICE_X21Y132_AO5),
.O6(CLBLM_R_X15Y132_SLICE_X21Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y116_SLICE_X0Y116_A5Q),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_BQ),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_B5Q),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X1Y115_A5Q),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X2Y115_A5Q),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_AQ),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X3Y115_A5Q),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X4Y115_A5Q),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(1'b0),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X16Y118_SLICE_X23Y118_AQ),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X15Y104_SLICE_X21Y104_BQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X16Y110_SLICE_X22Y110_AQ),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X15Y105_SLICE_X21Y105_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y141_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y141_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y142_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y142_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y143_IOB_X0Y143_IBUF (
.I(LIOB33_X0Y143_IOB_X0Y143_IPAD),
.O(LIOB33_X0Y143_IOB_X0Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y145_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y145_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y146_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y146_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y147_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y147_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y148_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y148_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y178_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y178_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y179_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y179_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y180_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y180_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y181_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y181_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y182_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y182_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y183_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y183_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y184_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y184_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y185_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y185_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y186_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y186_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y187_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y187_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y188_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y188_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y189_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y189_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y190_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y190_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y191_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y191_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y192_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y192_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y193_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y193_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y194_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y194_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y195_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y195_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y196_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y196_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y197_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y197_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y198_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y198_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y116_SLICE_X0Y116_AQ),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y149_IOB_X0Y149_IBUF (
.I(LIOB33_SING_X0Y149_IOB_X0Y149_IPAD),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y101_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.O(RIOB33_X105Y101_IOB_X1Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y102_OBUF (
.I(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.O(RIOB33_X105Y101_IOB_X1Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y103_OBUF (
.I(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.O(RIOB33_X105Y103_IOB_X1Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y104_OBUF (
.I(CLBLM_R_X11Y118_SLICE_X14Y118_A5Q),
.O(RIOB33_X105Y103_IOB_X1Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y105_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.O(RIOB33_X105Y105_IOB_X1Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y106_OBUF (
.I(CLBLM_L_X10Y119_SLICE_X13Y119_A5Q),
.O(RIOB33_X105Y105_IOB_X1Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUF (
.I(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUF (
.I(CLBLM_R_X11Y116_SLICE_X14Y116_A5Q),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X10Y116_B5Q),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y114_OBUF (
.I(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.O(RIOB33_X105Y113_IOB_X1Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(CLBLM_R_X15Y114_SLICE_X21Y114_AQ),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(CLBLM_L_X16Y114_SLICE_X22Y114_AQ),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(CLBLM_L_X16Y114_SLICE_X23Y114_BQ),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLM_L_X16Y116_SLICE_X23Y116_AQ),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLM_L_X16Y116_SLICE_X23Y116_BQ),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_R_X15Y116_SLICE_X20Y116_AQ),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLM_R_X15Y116_SLICE_X20Y116_BQ),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLM_R_X15Y115_SLICE_X20Y115_AQ),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLM_R_X15Y115_SLICE_X21Y115_AQ),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLM_L_X16Y115_SLICE_X22Y115_AQ),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_L_X16Y115_SLICE_X23Y115_AQ),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLM_L_X16Y115_SLICE_X23Y115_BQ),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_L_X16Y114_SLICE_X23Y114_AQ),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_R_X15Y114_SLICE_X20Y114_AQ),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_R_X15Y116_SLICE_X21Y116_AQ),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_R_X15Y116_SLICE_X21Y116_BQ),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_L_X16Y117_SLICE_X22Y117_AQ),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_L_X16Y117_SLICE_X22Y117_BQ),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_R_X15Y117_SLICE_X21Y117_BQ),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_L_X16Y118_SLICE_X23Y118_AQ),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_R_X15Y117_SLICE_X21Y117_AQ),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_R_X15Y117_SLICE_X20Y117_AQ),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLM_R_X15Y118_SLICE_X20Y118_AQ),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLM_R_X15Y119_SLICE_X20Y119_AQ),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_L_X16Y119_SLICE_X23Y119_AQ),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_L_X16Y119_SLICE_X22Y119_AQ),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_R_X15Y119_SLICE_X21Y119_AQ),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLM_R_X15Y119_SLICE_X21Y119_BQ),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLM_R_X15Y118_SLICE_X21Y118_AQ),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLM_R_X15Y132_SLICE_X21Y132_AQ),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLM_R_X15Y132_SLICE_X21Y132_BQ),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_R_X15Y132_SLICE_X21Y132_CQ),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_OBUF (
.I(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLM_R_X15Y132_SLICE_X21Y132_DQ),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_BMUX = CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_CMUX = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_AMUX = CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_AMUX = CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_CMUX = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_BMUX = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_AMUX = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AMUX = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_CMUX = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CMUX = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_BMUX = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CMUX = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CMUX = CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D = CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A = CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D = CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_AMUX = CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_BMUX = CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_AMUX = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_BMUX = CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_AMUX = CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_AMUX = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_BMUX = CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_CMUX = CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_DMUX = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_CMUX = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_DMUX = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_AMUX = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_AMUX = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_AMUX = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_BMUX = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_BMUX = CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_AMUX = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_AMUX = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_BMUX = CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_BMUX = CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_AMUX = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_BMUX = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CMUX = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_AMUX = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_AMUX = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CMUX = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AMUX = CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_DMUX = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_BMUX = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_DMUX = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_AMUX = CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_BMUX = CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A = CLBLM_L_X10Y100_SLICE_X12Y100_AO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B = CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C = CLBLM_L_X10Y100_SLICE_X12Y100_CO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D = CLBLM_L_X10Y100_SLICE_X12Y100_DO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_AMUX = CLBLM_L_X10Y100_SLICE_X12Y100_AO5;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A = CLBLM_L_X10Y100_SLICE_X13Y100_AO6;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B = CLBLM_L_X10Y100_SLICE_X13Y100_BO6;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C = CLBLM_L_X10Y100_SLICE_X13Y100_CO6;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D = CLBLM_L_X10Y100_SLICE_X13Y100_DO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A = CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C = CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D = CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_AMUX = CLBLM_L_X10Y101_SLICE_X12Y101_AO5;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B = CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C = CLBLM_L_X10Y101_SLICE_X13Y101_CO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D = CLBLM_L_X10Y101_SLICE_X13Y101_DO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_AMUX = CLBLM_L_X10Y101_SLICE_X13Y101_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_AMUX = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_AMUX = CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_BMUX = CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_AMUX = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_AMUX = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_BMUX = CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_AMUX = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_DMUX = CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_AMUX = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_AMUX = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_AMUX = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AMUX = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CMUX = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_AMUX = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_DMUX = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CMUX = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_DMUX = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_AMUX = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CMUX = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_AMUX = CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_AMUX = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_AMUX = CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CMUX = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CMUX = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_AMUX = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_BMUX = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CMUX = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_DMUX = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_AMUX = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_AMUX = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_AMUX = CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CMUX = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_AMUX = CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_AMUX = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CMUX = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_BMUX = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CMUX = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_BMUX = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CMUX = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_BMUX = CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_BMUX = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CMUX = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_BMUX = CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_BMUX = CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CMUX = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_CMUX = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_BMUX = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A = CLBLM_L_X12Y100_SLICE_X16Y100_AO6;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B = CLBLM_L_X12Y100_SLICE_X16Y100_BO6;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C = CLBLM_L_X12Y100_SLICE_X16Y100_CO6;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D = CLBLM_L_X12Y100_SLICE_X16Y100_DO6;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A = CLBLM_L_X12Y100_SLICE_X17Y100_AO6;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B = CLBLM_L_X12Y100_SLICE_X17Y100_BO6;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C = CLBLM_L_X12Y100_SLICE_X17Y100_CO6;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D = CLBLM_L_X12Y100_SLICE_X17Y100_DO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A = CLBLM_L_X12Y101_SLICE_X16Y101_AO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B = CLBLM_L_X12Y101_SLICE_X16Y101_BO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C = CLBLM_L_X12Y101_SLICE_X16Y101_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D = CLBLM_L_X12Y101_SLICE_X16Y101_DO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_AMUX = CLBLM_L_X12Y101_SLICE_X16Y101_AO5;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A = CLBLM_L_X12Y101_SLICE_X17Y101_AO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B = CLBLM_L_X12Y101_SLICE_X17Y101_BO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C = CLBLM_L_X12Y101_SLICE_X17Y101_CO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D = CLBLM_L_X12Y101_SLICE_X17Y101_DO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_CMUX = CLBLM_L_X12Y101_SLICE_X17Y101_CO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_DMUX = CLBLM_L_X12Y101_SLICE_X17Y101_DO5;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A = CLBLM_L_X12Y102_SLICE_X16Y102_AO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B = CLBLM_L_X12Y102_SLICE_X16Y102_BO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C = CLBLM_L_X12Y102_SLICE_X16Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D = CLBLM_L_X12Y102_SLICE_X16Y102_DO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_CMUX = CLBLM_L_X12Y102_SLICE_X16Y102_CO5;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A = CLBLM_L_X12Y102_SLICE_X17Y102_AO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B = CLBLM_L_X12Y102_SLICE_X17Y102_BO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C = CLBLM_L_X12Y102_SLICE_X17Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D = CLBLM_L_X12Y102_SLICE_X17Y102_DO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_AMUX = CLBLM_L_X12Y102_SLICE_X17Y102_AO5;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A = CLBLM_L_X12Y103_SLICE_X16Y103_AO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B = CLBLM_L_X12Y103_SLICE_X16Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C = CLBLM_L_X12Y103_SLICE_X16Y103_CO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D = CLBLM_L_X12Y103_SLICE_X16Y103_DO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_BMUX = CLBLM_L_X12Y103_SLICE_X16Y103_BO5;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A = CLBLM_L_X12Y103_SLICE_X17Y103_AO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B = CLBLM_L_X12Y103_SLICE_X17Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C = CLBLM_L_X12Y103_SLICE_X17Y103_CO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D = CLBLM_L_X12Y103_SLICE_X17Y103_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_CMUX = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A = CLBLM_L_X12Y104_SLICE_X17Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B = CLBLM_L_X12Y104_SLICE_X17Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C = CLBLM_L_X12Y104_SLICE_X17Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D = CLBLM_L_X12Y104_SLICE_X17Y104_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_DMUX = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_AMUX = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_AMUX = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_AMUX = CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_AMUX = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_DMUX = CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_CMUX = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_BMUX = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_AMUX = CLBLM_L_X12Y111_SLICE_X16Y111_AO5;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A = CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B = CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C = CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D = CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B = CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C = CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D = CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A = CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C = CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_BMUX = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_DMUX = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_AMUX = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_BMUX = CLBLM_L_X12Y113_SLICE_X16Y113_BO5;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_CMUX = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A = CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B = CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C = CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_AMUX = CLBLM_L_X12Y113_SLICE_X17Y113_AO5;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A = CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A = CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B = CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C = CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D = CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_AMUX = CLBLM_L_X12Y115_SLICE_X16Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_BMUX = CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CMUX = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_AMUX = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_BMUX = CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A = CLBLM_L_X12Y116_SLICE_X16Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_AMUX = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_BMUX = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CMUX = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A = CLBLM_L_X12Y116_SLICE_X17Y116_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B = CLBLM_L_X12Y116_SLICE_X17Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_AMUX = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_BMUX = CLBLM_L_X12Y116_SLICE_X17Y116_BO5;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_CMUX = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_AMUX = CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_BMUX = CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A = CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D = CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A = CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_DMUX = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A = CLBLM_L_X12Y122_SLICE_X16Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A = CLBLM_L_X12Y122_SLICE_X17Y122_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_DMUX = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A = CLBLM_L_X12Y123_SLICE_X16Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B = CLBLM_L_X12Y123_SLICE_X16Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_CMUX = CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A = CLBLM_L_X12Y123_SLICE_X17Y123_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A = CLBLM_L_X12Y124_SLICE_X16Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A = CLBLM_L_X12Y124_SLICE_X17Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_DMUX = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A = CLBLM_L_X12Y125_SLICE_X16Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B = CLBLM_L_X12Y125_SLICE_X16Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_DMUX = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_BMUX = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A = CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CMUX = CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_CMUX = CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A = CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_BMUX = CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_AMUX = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_BMUX = CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_BMUX = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A = CLBLM_L_X16Y101_SLICE_X22Y101_AO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B = CLBLM_L_X16Y101_SLICE_X22Y101_BO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C = CLBLM_L_X16Y101_SLICE_X22Y101_CO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D = CLBLM_L_X16Y101_SLICE_X22Y101_DO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_BMUX = CLBLM_L_X16Y101_SLICE_X22Y101_BO5;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A = CLBLM_L_X16Y101_SLICE_X23Y101_AO6;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B = CLBLM_L_X16Y101_SLICE_X23Y101_BO6;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C = CLBLM_L_X16Y101_SLICE_X23Y101_CO6;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D = CLBLM_L_X16Y101_SLICE_X23Y101_DO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A = CLBLM_L_X16Y102_SLICE_X22Y102_AO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B = CLBLM_L_X16Y102_SLICE_X22Y102_BO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C = CLBLM_L_X16Y102_SLICE_X22Y102_CO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D = CLBLM_L_X16Y102_SLICE_X22Y102_DO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_BMUX = CLBLM_L_X16Y102_SLICE_X22Y102_BO5;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_CMUX = CLBLM_L_X16Y102_SLICE_X22Y102_CO5;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A = CLBLM_L_X16Y102_SLICE_X23Y102_AO6;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B = CLBLM_L_X16Y102_SLICE_X23Y102_BO6;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C = CLBLM_L_X16Y102_SLICE_X23Y102_CO6;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D = CLBLM_L_X16Y102_SLICE_X23Y102_DO6;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_AMUX = CLBLM_L_X16Y102_SLICE_X23Y102_AO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A = CLBLM_L_X16Y103_SLICE_X22Y103_AO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B = CLBLM_L_X16Y103_SLICE_X22Y103_BO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C = CLBLM_L_X16Y103_SLICE_X22Y103_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D = CLBLM_L_X16Y103_SLICE_X22Y103_DO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_DMUX = CLBLM_L_X16Y103_SLICE_X22Y103_DO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A = CLBLM_L_X16Y103_SLICE_X23Y103_AO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B = CLBLM_L_X16Y103_SLICE_X23Y103_BO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D = CLBLM_L_X16Y103_SLICE_X23Y103_DO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A = CLBLM_L_X16Y104_SLICE_X22Y104_AO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B = CLBLM_L_X16Y104_SLICE_X22Y104_BO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C = CLBLM_L_X16Y104_SLICE_X22Y104_CO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D = CLBLM_L_X16Y104_SLICE_X22Y104_DO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A = CLBLM_L_X16Y104_SLICE_X23Y104_AO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B = CLBLM_L_X16Y104_SLICE_X23Y104_BO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C = CLBLM_L_X16Y104_SLICE_X23Y104_CO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D = CLBLM_L_X16Y104_SLICE_X23Y104_DO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A = CLBLM_L_X16Y105_SLICE_X22Y105_AO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B = CLBLM_L_X16Y105_SLICE_X22Y105_BO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C = CLBLM_L_X16Y105_SLICE_X22Y105_CO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D = CLBLM_L_X16Y105_SLICE_X22Y105_DO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A = CLBLM_L_X16Y105_SLICE_X23Y105_AO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B = CLBLM_L_X16Y105_SLICE_X23Y105_BO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C = CLBLM_L_X16Y105_SLICE_X23Y105_CO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D = CLBLM_L_X16Y105_SLICE_X23Y105_DO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_AMUX = CLBLM_L_X16Y105_SLICE_X23Y105_AO5;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A = CLBLM_L_X16Y106_SLICE_X22Y106_AO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B = CLBLM_L_X16Y106_SLICE_X22Y106_BO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C = CLBLM_L_X16Y106_SLICE_X22Y106_CO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D = CLBLM_L_X16Y106_SLICE_X22Y106_DO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_BMUX = CLBLM_L_X16Y106_SLICE_X22Y106_BO5;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_CMUX = CLBLM_L_X16Y106_SLICE_X22Y106_CO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A = CLBLM_L_X16Y106_SLICE_X23Y106_AO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B = CLBLM_L_X16Y106_SLICE_X23Y106_BO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C = CLBLM_L_X16Y106_SLICE_X23Y106_CO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D = CLBLM_L_X16Y106_SLICE_X23Y106_DO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_AMUX = CLBLM_L_X16Y106_SLICE_X23Y106_AO5;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_BMUX = CLBLM_L_X16Y106_SLICE_X23Y106_BO5;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_CMUX = CLBLM_L_X16Y106_SLICE_X23Y106_CO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A = CLBLM_L_X16Y107_SLICE_X22Y107_AO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B = CLBLM_L_X16Y107_SLICE_X22Y107_BO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C = CLBLM_L_X16Y107_SLICE_X22Y107_CO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D = CLBLM_L_X16Y107_SLICE_X22Y107_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A = CLBLM_L_X16Y107_SLICE_X23Y107_AO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B = CLBLM_L_X16Y107_SLICE_X23Y107_BO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C = CLBLM_L_X16Y107_SLICE_X23Y107_CO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D = CLBLM_L_X16Y107_SLICE_X23Y107_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_DMUX = CLBLM_L_X16Y107_SLICE_X23Y107_DO5;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A = CLBLM_L_X16Y108_SLICE_X22Y108_AO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B = CLBLM_L_X16Y108_SLICE_X22Y108_BO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C = CLBLM_L_X16Y108_SLICE_X22Y108_CO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D = CLBLM_L_X16Y108_SLICE_X22Y108_DO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_AMUX = CLBLM_L_X16Y108_SLICE_X22Y108_AO5;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A = CLBLM_L_X16Y108_SLICE_X23Y108_AO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B = CLBLM_L_X16Y108_SLICE_X23Y108_BO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C = CLBLM_L_X16Y108_SLICE_X23Y108_CO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D = CLBLM_L_X16Y108_SLICE_X23Y108_DO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A = CLBLM_L_X16Y109_SLICE_X22Y109_AO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B = CLBLM_L_X16Y109_SLICE_X22Y109_BO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C = CLBLM_L_X16Y109_SLICE_X22Y109_CO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D = CLBLM_L_X16Y109_SLICE_X22Y109_DO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_AMUX = CLBLM_L_X16Y109_SLICE_X22Y109_AO5;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_BMUX = CLBLM_L_X16Y109_SLICE_X22Y109_BO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A = CLBLM_L_X16Y109_SLICE_X23Y109_AO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B = CLBLM_L_X16Y109_SLICE_X23Y109_BO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C = CLBLM_L_X16Y109_SLICE_X23Y109_CO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D = CLBLM_L_X16Y109_SLICE_X23Y109_DO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_AMUX = CLBLM_L_X16Y109_SLICE_X23Y109_AO5;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A = CLBLM_L_X16Y110_SLICE_X22Y110_AO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B = CLBLM_L_X16Y110_SLICE_X22Y110_BO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C = CLBLM_L_X16Y110_SLICE_X22Y110_CO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D = CLBLM_L_X16Y110_SLICE_X22Y110_DO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A = CLBLM_L_X16Y110_SLICE_X23Y110_AO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B = CLBLM_L_X16Y110_SLICE_X23Y110_BO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C = CLBLM_L_X16Y110_SLICE_X23Y110_CO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D = CLBLM_L_X16Y110_SLICE_X23Y110_DO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_AMUX = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A = CLBLM_L_X16Y111_SLICE_X22Y111_AO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B = CLBLM_L_X16Y111_SLICE_X22Y111_BO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C = CLBLM_L_X16Y111_SLICE_X22Y111_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D = CLBLM_L_X16Y111_SLICE_X22Y111_DO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A = CLBLM_L_X16Y111_SLICE_X23Y111_AO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B = CLBLM_L_X16Y111_SLICE_X23Y111_BO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C = CLBLM_L_X16Y111_SLICE_X23Y111_CO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D = CLBLM_L_X16Y111_SLICE_X23Y111_DO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_BMUX = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A = CLBLM_L_X16Y113_SLICE_X22Y113_AO6;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B = CLBLM_L_X16Y113_SLICE_X22Y113_BO6;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C = CLBLM_L_X16Y113_SLICE_X22Y113_CO6;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D = CLBLM_L_X16Y113_SLICE_X22Y113_DO6;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_AMUX = CLBLM_L_X16Y113_SLICE_X22Y113_AO5;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_BMUX = CLBLM_L_X16Y113_SLICE_X22Y113_BO5;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_CMUX = CLBLM_L_X16Y113_SLICE_X22Y113_CO5;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A = CLBLM_L_X16Y113_SLICE_X23Y113_AO6;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B = CLBLM_L_X16Y113_SLICE_X23Y113_BO6;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C = CLBLM_L_X16Y113_SLICE_X23Y113_CO6;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D = CLBLM_L_X16Y113_SLICE_X23Y113_DO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A = CLBLM_L_X16Y114_SLICE_X22Y114_AO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B = CLBLM_L_X16Y114_SLICE_X22Y114_BO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C = CLBLM_L_X16Y114_SLICE_X22Y114_CO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D = CLBLM_L_X16Y114_SLICE_X22Y114_DO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_BMUX = CLBLM_L_X16Y114_SLICE_X22Y114_BO5;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_CMUX = CLBLM_L_X16Y114_SLICE_X22Y114_CO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A = CLBLM_L_X16Y114_SLICE_X23Y114_AO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B = CLBLM_L_X16Y114_SLICE_X23Y114_BO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C = CLBLM_L_X16Y114_SLICE_X23Y114_CO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D = CLBLM_L_X16Y114_SLICE_X23Y114_DO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A = CLBLM_L_X16Y115_SLICE_X22Y115_AO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B = CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C = CLBLM_L_X16Y115_SLICE_X22Y115_CO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D = CLBLM_L_X16Y115_SLICE_X22Y115_DO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A = CLBLM_L_X16Y115_SLICE_X23Y115_AO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B = CLBLM_L_X16Y115_SLICE_X23Y115_BO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C = CLBLM_L_X16Y115_SLICE_X23Y115_CO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D = CLBLM_L_X16Y115_SLICE_X23Y115_DO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_CMUX = CLBLM_L_X16Y115_SLICE_X23Y115_CO5;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A = CLBLM_L_X16Y116_SLICE_X22Y116_AO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B = CLBLM_L_X16Y116_SLICE_X22Y116_BO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C = CLBLM_L_X16Y116_SLICE_X22Y116_CO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D = CLBLM_L_X16Y116_SLICE_X22Y116_DO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_AMUX = CLBLM_L_X16Y116_SLICE_X22Y116_AO5;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_BMUX = CLBLM_L_X16Y116_SLICE_X22Y116_BO5;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_CMUX = CLBLM_L_X16Y116_SLICE_X22Y116_CO5;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A = CLBLM_L_X16Y116_SLICE_X23Y116_AO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B = CLBLM_L_X16Y116_SLICE_X23Y116_BO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C = CLBLM_L_X16Y116_SLICE_X23Y116_CO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D = CLBLM_L_X16Y116_SLICE_X23Y116_DO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A = CLBLM_L_X16Y117_SLICE_X22Y117_AO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B = CLBLM_L_X16Y117_SLICE_X22Y117_BO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C = CLBLM_L_X16Y117_SLICE_X22Y117_CO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D = CLBLM_L_X16Y117_SLICE_X22Y117_DO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A = CLBLM_L_X16Y117_SLICE_X23Y117_AO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B = CLBLM_L_X16Y117_SLICE_X23Y117_BO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C = CLBLM_L_X16Y117_SLICE_X23Y117_CO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D = CLBLM_L_X16Y117_SLICE_X23Y117_DO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_AMUX = CLBLM_L_X16Y117_SLICE_X23Y117_AO5;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A = CLBLM_L_X16Y118_SLICE_X22Y118_AO6;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B = CLBLM_L_X16Y118_SLICE_X22Y118_BO6;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C = CLBLM_L_X16Y118_SLICE_X22Y118_CO6;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D = CLBLM_L_X16Y118_SLICE_X22Y118_DO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A = CLBLM_L_X16Y118_SLICE_X23Y118_AO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B = CLBLM_L_X16Y118_SLICE_X23Y118_BO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C = CLBLM_L_X16Y118_SLICE_X23Y118_CO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D = CLBLM_L_X16Y118_SLICE_X23Y118_DO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A = CLBLM_L_X16Y119_SLICE_X22Y119_AO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B = CLBLM_L_X16Y119_SLICE_X22Y119_BO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C = CLBLM_L_X16Y119_SLICE_X22Y119_CO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D = CLBLM_L_X16Y119_SLICE_X22Y119_DO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_BMUX = CLBLM_L_X16Y119_SLICE_X22Y119_BO5;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_CMUX = CLBLM_L_X16Y119_SLICE_X22Y119_CO5;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A = CLBLM_L_X16Y119_SLICE_X23Y119_AO6;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B = CLBLM_L_X16Y119_SLICE_X23Y119_BO6;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C = CLBLM_L_X16Y119_SLICE_X23Y119_CO6;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D = CLBLM_L_X16Y119_SLICE_X23Y119_DO6;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A = CLBLM_L_X16Y121_SLICE_X22Y121_AO6;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B = CLBLM_L_X16Y121_SLICE_X22Y121_BO6;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C = CLBLM_L_X16Y121_SLICE_X22Y121_CO6;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D = CLBLM_L_X16Y121_SLICE_X22Y121_DO6;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A = CLBLM_L_X16Y121_SLICE_X23Y121_AO6;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B = CLBLM_L_X16Y121_SLICE_X23Y121_BO6;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C = CLBLM_L_X16Y121_SLICE_X23Y121_CO6;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D = CLBLM_L_X16Y121_SLICE_X23Y121_DO6;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A = CLBLM_L_X16Y123_SLICE_X22Y123_AO6;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C = CLBLM_L_X16Y123_SLICE_X22Y123_CO6;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D = CLBLM_L_X16Y123_SLICE_X22Y123_DO6;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_AMUX = CLBLM_L_X16Y123_SLICE_X22Y123_AO5;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A = CLBLM_L_X16Y123_SLICE_X23Y123_AO6;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B = CLBLM_L_X16Y123_SLICE_X23Y123_BO6;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C = CLBLM_L_X16Y123_SLICE_X23Y123_CO6;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D = CLBLM_L_X16Y123_SLICE_X23Y123_DO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A = CLBLM_L_X16Y125_SLICE_X22Y125_AO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B = CLBLM_L_X16Y125_SLICE_X22Y125_BO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C = CLBLM_L_X16Y125_SLICE_X22Y125_CO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_BMUX = CLBLM_L_X16Y125_SLICE_X22Y125_BO5;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_CMUX = CLBLM_L_X16Y125_SLICE_X22Y125_CO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A = CLBLM_L_X16Y125_SLICE_X23Y125_AO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D = CLBLM_L_X16Y125_SLICE_X23Y125_DO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_AMUX = CLBLM_L_X16Y125_SLICE_X23Y125_AO5;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A = CLBLM_L_X16Y126_SLICE_X22Y126_AO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B = CLBLM_L_X16Y126_SLICE_X22Y126_BO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C = CLBLM_L_X16Y126_SLICE_X22Y126_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D = CLBLM_L_X16Y126_SLICE_X22Y126_DO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_BMUX = CLBLM_L_X16Y126_SLICE_X22Y126_BO5;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D = CLBLM_L_X16Y126_SLICE_X23Y126_DO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_AMUX = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_BMUX = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_AMUX = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_BMUX = CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AMUX = CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CMUX = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CMUX = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_BMUX = CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_BMUX = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_DMUX = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_AMUX = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_AMUX = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_AMUX = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_BMUX = CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_DMUX = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_BMUX = CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_CMUX = CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_AMUX = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_AMUX = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_CMUX = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CMUX = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CMUX = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_BMUX = CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_BMUX = CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_BMUX = CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_BMUX = CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_DMUX = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_BMUX = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CMUX = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_BMUX = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_AMUX = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_BMUX = CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_AMUX = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_BMUX = CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_AMUX = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_AMUX = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_CMUX = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_AMUX = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_AMUX = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_AMUX = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_CMUX = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_BMUX = CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_CMUX = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CMUX = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_BMUX = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_CMUX = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_AMUX = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_BMUX = CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_CMUX = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_AMUX = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CMUX = CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_DMUX = CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_AMUX = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CMUX = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_AMUX = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_BMUX = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_AMUX = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_BMUX = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CMUX = CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_AMUX = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CMUX = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CMUX = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_BMUX = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_AMUX = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_BMUX = CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CMUX = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_BMUX = CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CMUX = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_BMUX = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CMUX = CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_AMUX = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_AMUX = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_BMUX = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CMUX = CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_AMUX = CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_AMUX = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A = CLBLM_R_X11Y100_SLICE_X14Y100_AO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C = CLBLM_R_X11Y100_SLICE_X14Y100_CO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D = CLBLM_R_X11Y100_SLICE_X14Y100_DO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_AMUX = CLBLM_R_X11Y100_SLICE_X14Y100_AO5;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A = CLBLM_R_X11Y100_SLICE_X15Y100_AO6;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B = CLBLM_R_X11Y100_SLICE_X15Y100_BO6;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C = CLBLM_R_X11Y100_SLICE_X15Y100_CO6;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D = CLBLM_R_X11Y100_SLICE_X15Y100_DO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A = CLBLM_R_X11Y101_SLICE_X14Y101_AO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B = CLBLM_R_X11Y101_SLICE_X14Y101_BO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C = CLBLM_R_X11Y101_SLICE_X14Y101_CO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D = CLBLM_R_X11Y101_SLICE_X14Y101_DO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A = CLBLM_R_X11Y101_SLICE_X15Y101_AO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B = CLBLM_R_X11Y101_SLICE_X15Y101_BO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C = CLBLM_R_X11Y101_SLICE_X15Y101_CO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D = CLBLM_R_X11Y101_SLICE_X15Y101_DO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_AMUX = CLBLM_R_X11Y101_SLICE_X15Y101_AO5;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A = CLBLM_R_X11Y102_SLICE_X14Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B = CLBLM_R_X11Y102_SLICE_X14Y102_BO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C = CLBLM_R_X11Y102_SLICE_X14Y102_CO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D = CLBLM_R_X11Y102_SLICE_X14Y102_DO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_AMUX = CLBLM_R_X11Y102_SLICE_X14Y102_AO5;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A = CLBLM_R_X11Y102_SLICE_X15Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B = CLBLM_R_X11Y102_SLICE_X15Y102_BO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C = CLBLM_R_X11Y102_SLICE_X15Y102_CO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D = CLBLM_R_X11Y102_SLICE_X15Y102_DO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_AMUX = CLBLM_R_X11Y102_SLICE_X15Y102_AO5;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_CMUX = CLBLM_R_X11Y102_SLICE_X15Y102_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B = CLBLM_R_X11Y103_SLICE_X14Y103_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C = CLBLM_R_X11Y103_SLICE_X14Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D = CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_CMUX = CLBLM_R_X11Y103_SLICE_X14Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_DMUX = CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A = CLBLM_R_X11Y103_SLICE_X15Y103_AO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B = CLBLM_R_X11Y103_SLICE_X15Y103_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C = CLBLM_R_X11Y103_SLICE_X15Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D = CLBLM_R_X11Y103_SLICE_X15Y103_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_CMUX = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_AMUX = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_DMUX = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_DMUX = CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_AMUX = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_CMUX = CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_CMUX = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_BMUX = CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_BMUX = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_BMUX = CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_CMUX = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_AMUX = CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_BMUX = CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_CMUX = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_AMUX = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_BMUX = CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_CMUX = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_AMUX = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_AMUX = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_CMUX = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_AMUX = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_BMUX = CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_AMUX = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CMUX = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CMUX = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_AMUX = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_AMUX = CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CMUX = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A = CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B = CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_AMUX = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A = CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_BMUX = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_BMUX = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_AMUX = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_BMUX = CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CMUX = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_AMUX = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_AMUX = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_BMUX = CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_CMUX = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_DMUX = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_AMUX = CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_CMUX = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_BMUX = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A = CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A = CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_AMUX = CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_BMUX = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_BMUX = CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_BMUX = CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CMUX = CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A = CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CMUX = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A = CLBLM_R_X13Y100_SLICE_X18Y100_AO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B = CLBLM_R_X13Y100_SLICE_X18Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C = CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D = CLBLM_R_X13Y100_SLICE_X18Y100_DO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_BMUX = CLBLM_R_X13Y100_SLICE_X18Y100_BO5;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_DMUX = CLBLM_R_X13Y100_SLICE_X18Y100_DO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B = CLBLM_R_X13Y100_SLICE_X19Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C = CLBLM_R_X13Y100_SLICE_X19Y100_CO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D = CLBLM_R_X13Y100_SLICE_X19Y100_DO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_BMUX = CLBLM_R_X13Y100_SLICE_X19Y100_BO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A = CLBLM_R_X13Y101_SLICE_X18Y101_AO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B = CLBLM_R_X13Y101_SLICE_X18Y101_BO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C = CLBLM_R_X13Y101_SLICE_X18Y101_CO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D = CLBLM_R_X13Y101_SLICE_X18Y101_DO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_BMUX = CLBLM_R_X13Y101_SLICE_X18Y101_BO5;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A = CLBLM_R_X13Y101_SLICE_X19Y101_AO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B = CLBLM_R_X13Y101_SLICE_X19Y101_BO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C = CLBLM_R_X13Y101_SLICE_X19Y101_CO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_AMUX = CLBLM_R_X13Y101_SLICE_X19Y101_AO5;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A = CLBLM_R_X13Y102_SLICE_X18Y102_AO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B = CLBLM_R_X13Y102_SLICE_X18Y102_BO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C = CLBLM_R_X13Y102_SLICE_X18Y102_CO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D = CLBLM_R_X13Y102_SLICE_X18Y102_DO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_CMUX = CLBLM_R_X13Y102_SLICE_X18Y102_CO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A = CLBLM_R_X13Y102_SLICE_X19Y102_AO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B = CLBLM_R_X13Y102_SLICE_X19Y102_BO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C = CLBLM_R_X13Y102_SLICE_X19Y102_CO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D = CLBLM_R_X13Y102_SLICE_X19Y102_DO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_AMUX = CLBLM_R_X13Y102_SLICE_X19Y102_AO5;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A = CLBLM_R_X13Y103_SLICE_X18Y103_AO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B = CLBLM_R_X13Y103_SLICE_X18Y103_BO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C = CLBLM_R_X13Y103_SLICE_X18Y103_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D = CLBLM_R_X13Y103_SLICE_X18Y103_DO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_BMUX = CLBLM_R_X13Y103_SLICE_X18Y103_BO5;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A = CLBLM_R_X13Y103_SLICE_X19Y103_AO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B = CLBLM_R_X13Y103_SLICE_X19Y103_BO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C = CLBLM_R_X13Y103_SLICE_X19Y103_CO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D = CLBLM_R_X13Y103_SLICE_X19Y103_DO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_AMUX = CLBLM_R_X13Y103_SLICE_X19Y103_AO5;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A = CLBLM_R_X13Y104_SLICE_X18Y104_AO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B = CLBLM_R_X13Y104_SLICE_X18Y104_BO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C = CLBLM_R_X13Y104_SLICE_X18Y104_CO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D = CLBLM_R_X13Y104_SLICE_X18Y104_DO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A = CLBLM_R_X13Y104_SLICE_X19Y104_AO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B = CLBLM_R_X13Y104_SLICE_X19Y104_BO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C = CLBLM_R_X13Y104_SLICE_X19Y104_CO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D = CLBLM_R_X13Y104_SLICE_X19Y104_DO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_AMUX = CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A = CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D = CLBLM_R_X13Y106_SLICE_X19Y106_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D = CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_AMUX = CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A = CLBLM_R_X13Y107_SLICE_X19Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B = CLBLM_R_X13Y107_SLICE_X19Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C = CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D = CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C = CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D = CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_AMUX = CLBLM_R_X13Y108_SLICE_X19Y108_AO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_DMUX = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B = CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C = CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D = CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A = CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B = CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C = CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D = CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A = CLBLM_R_X13Y111_SLICE_X18Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B = CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_BMUX = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_DMUX = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B = CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C = CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D = CLBLM_R_X13Y111_SLICE_X19Y111_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B = CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_AMUX = CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_BMUX = CLBLM_R_X13Y112_SLICE_X18Y112_BO5;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B = CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_CMUX = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A = CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B = CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C = CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A = CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_AMUX = CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A = CLBLM_R_X13Y114_SLICE_X18Y114_AO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B = CLBLM_R_X13Y114_SLICE_X18Y114_BO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C = CLBLM_R_X13Y114_SLICE_X18Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D = CLBLM_R_X13Y114_SLICE_X18Y114_DO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_AMUX = CLBLM_R_X13Y114_SLICE_X18Y114_AO5;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A = CLBLM_R_X13Y114_SLICE_X19Y114_AO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C = CLBLM_R_X13Y114_SLICE_X19Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D = CLBLM_R_X13Y114_SLICE_X19Y114_DO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_AMUX = CLBLM_R_X13Y114_SLICE_X19Y114_AO5;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A = CLBLM_R_X13Y115_SLICE_X18Y115_AO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B = CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D = CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_AMUX = CLBLM_R_X13Y115_SLICE_X18Y115_AO5;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A = CLBLM_R_X13Y115_SLICE_X19Y115_AO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B = CLBLM_R_X13Y115_SLICE_X19Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C = CLBLM_R_X13Y115_SLICE_X19Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D = CLBLM_R_X13Y115_SLICE_X19Y115_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B = CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A = CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B = CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C = CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D = CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B = CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C = CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D = CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_AMUX = CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A = CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B = CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C = CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D = CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A = CLBLM_R_X13Y119_SLICE_X18Y119_AO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C = CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_BMUX = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A = CLBLM_R_X13Y119_SLICE_X19Y119_AO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B = CLBLM_R_X13Y119_SLICE_X19Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C = CLBLM_R_X13Y119_SLICE_X19Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D = CLBLM_R_X13Y119_SLICE_X19Y119_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A = CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A = CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C = CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_CMUX = CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A = CLBLM_R_X13Y121_SLICE_X18Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B = CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A = CLBLM_R_X13Y121_SLICE_X19Y121_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B = CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C = CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A = CLBLM_R_X13Y122_SLICE_X18Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B = CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A = CLBLM_R_X13Y122_SLICE_X19Y122_AO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A = CLBLM_R_X13Y123_SLICE_X18Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B = CLBLM_R_X13Y123_SLICE_X18Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A = CLBLM_R_X13Y123_SLICE_X19Y123_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B = CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C = CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A = CLBLM_R_X13Y124_SLICE_X18Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B = CLBLM_R_X13Y124_SLICE_X18Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A = CLBLM_R_X13Y124_SLICE_X19Y124_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B = CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D = CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_BMUX = CLBLM_R_X13Y124_SLICE_X19Y124_BO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A = CLBLM_R_X13Y125_SLICE_X18Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D = CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_BMUX = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A = CLBLM_R_X13Y125_SLICE_X19Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D = CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A = CLBLM_R_X13Y126_SLICE_X18Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B = CLBLM_R_X13Y126_SLICE_X18Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A = CLBLM_R_X13Y126_SLICE_X19Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B = CLBLM_R_X13Y126_SLICE_X19Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D = CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_AMUX = CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CMUX = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A = CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_BMUX = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_AMUX = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_AMUX = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D = CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_AMUX = CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_BMUX = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A = CLBLM_R_X15Y100_SLICE_X20Y100_AO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B = CLBLM_R_X15Y100_SLICE_X20Y100_BO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C = CLBLM_R_X15Y100_SLICE_X20Y100_CO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D = CLBLM_R_X15Y100_SLICE_X20Y100_DO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_BMUX = CLBLM_R_X15Y100_SLICE_X20Y100_BO5;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_DMUX = CLBLM_R_X15Y100_SLICE_X20Y100_DO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A = CLBLM_R_X15Y100_SLICE_X21Y100_AO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B = CLBLM_R_X15Y100_SLICE_X21Y100_BO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C = CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D = CLBLM_R_X15Y100_SLICE_X21Y100_DO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A = CLBLM_R_X15Y101_SLICE_X20Y101_AO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B = CLBLM_R_X15Y101_SLICE_X20Y101_BO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C = CLBLM_R_X15Y101_SLICE_X20Y101_CO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D = CLBLM_R_X15Y101_SLICE_X20Y101_DO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_AMUX = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_BMUX = CLBLM_R_X15Y101_SLICE_X20Y101_BO5;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A = CLBLM_R_X15Y101_SLICE_X21Y101_AO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B = CLBLM_R_X15Y101_SLICE_X21Y101_BO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C = CLBLM_R_X15Y101_SLICE_X21Y101_CO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D = CLBLM_R_X15Y101_SLICE_X21Y101_DO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_AMUX = CLBLM_R_X15Y101_SLICE_X21Y101_AO5;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_BMUX = CLBLM_R_X15Y101_SLICE_X21Y101_BO5;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A = CLBLM_R_X15Y102_SLICE_X20Y102_AO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B = CLBLM_R_X15Y102_SLICE_X20Y102_BO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C = CLBLM_R_X15Y102_SLICE_X20Y102_CO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D = CLBLM_R_X15Y102_SLICE_X20Y102_DO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A = CLBLM_R_X15Y102_SLICE_X21Y102_AO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B = CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C = CLBLM_R_X15Y102_SLICE_X21Y102_CO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D = CLBLM_R_X15Y102_SLICE_X21Y102_DO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_AMUX = CLBLM_R_X15Y102_SLICE_X21Y102_AO5;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A = CLBLM_R_X15Y103_SLICE_X20Y103_AO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B = CLBLM_R_X15Y103_SLICE_X20Y103_BO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C = CLBLM_R_X15Y103_SLICE_X20Y103_CO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D = CLBLM_R_X15Y103_SLICE_X20Y103_DO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_AMUX = CLBLM_R_X15Y103_SLICE_X20Y103_AO5;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_CMUX = CLBLM_R_X15Y103_SLICE_X20Y103_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A = CLBLM_R_X15Y103_SLICE_X21Y103_AO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B = CLBLM_R_X15Y103_SLICE_X21Y103_BO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C = CLBLM_R_X15Y103_SLICE_X21Y103_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D = CLBLM_R_X15Y103_SLICE_X21Y103_DO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_AMUX = CLBLM_R_X15Y103_SLICE_X21Y103_AO5;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A = CLBLM_R_X15Y104_SLICE_X20Y104_AO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B = CLBLM_R_X15Y104_SLICE_X20Y104_BO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C = CLBLM_R_X15Y104_SLICE_X20Y104_CO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D = CLBLM_R_X15Y104_SLICE_X20Y104_DO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A = CLBLM_R_X15Y104_SLICE_X21Y104_AO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B = CLBLM_R_X15Y104_SLICE_X21Y104_BO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C = CLBLM_R_X15Y104_SLICE_X21Y104_CO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D = CLBLM_R_X15Y104_SLICE_X21Y104_DO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A = CLBLM_R_X15Y105_SLICE_X20Y105_AO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B = CLBLM_R_X15Y105_SLICE_X20Y105_BO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C = CLBLM_R_X15Y105_SLICE_X20Y105_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D = CLBLM_R_X15Y105_SLICE_X20Y105_DO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_DMUX = CLBLM_R_X15Y105_SLICE_X20Y105_DO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A = CLBLM_R_X15Y105_SLICE_X21Y105_AO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B = CLBLM_R_X15Y105_SLICE_X21Y105_BO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C = CLBLM_R_X15Y105_SLICE_X21Y105_CO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D = CLBLM_R_X15Y105_SLICE_X21Y105_DO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_BMUX = CLBLM_R_X15Y105_SLICE_X21Y105_BO5;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A = CLBLM_R_X15Y106_SLICE_X20Y106_AO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B = CLBLM_R_X15Y106_SLICE_X20Y106_BO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C = CLBLM_R_X15Y106_SLICE_X20Y106_CO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D = CLBLM_R_X15Y106_SLICE_X20Y106_DO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_DMUX = CLBLM_R_X15Y106_SLICE_X20Y106_DO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A = CLBLM_R_X15Y106_SLICE_X21Y106_AO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B = CLBLM_R_X15Y106_SLICE_X21Y106_BO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C = CLBLM_R_X15Y106_SLICE_X21Y106_CO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D = CLBLM_R_X15Y106_SLICE_X21Y106_DO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_BMUX = CLBLM_R_X15Y106_SLICE_X21Y106_BO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A = CLBLM_R_X15Y107_SLICE_X20Y107_AO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B = CLBLM_R_X15Y107_SLICE_X20Y107_BO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C = CLBLM_R_X15Y107_SLICE_X20Y107_CO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D = CLBLM_R_X15Y107_SLICE_X20Y107_DO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_BMUX = CLBLM_R_X15Y107_SLICE_X20Y107_BO5;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_CMUX = CLBLM_R_X15Y107_SLICE_X20Y107_CO5;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A = CLBLM_R_X15Y107_SLICE_X21Y107_AO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B = CLBLM_R_X15Y107_SLICE_X21Y107_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C = CLBLM_R_X15Y107_SLICE_X21Y107_CO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D = CLBLM_R_X15Y107_SLICE_X21Y107_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_AMUX = CLBLM_R_X15Y107_SLICE_X21Y107_AO5;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A = CLBLM_R_X15Y108_SLICE_X20Y108_AO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B = CLBLM_R_X15Y108_SLICE_X20Y108_BO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C = CLBLM_R_X15Y108_SLICE_X20Y108_CO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D = CLBLM_R_X15Y108_SLICE_X20Y108_DO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_AMUX = CLBLM_R_X15Y108_SLICE_X20Y108_AO5;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A = CLBLM_R_X15Y108_SLICE_X21Y108_AO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B = CLBLM_R_X15Y108_SLICE_X21Y108_BO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C = CLBLM_R_X15Y108_SLICE_X21Y108_CO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D = CLBLM_R_X15Y108_SLICE_X21Y108_DO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_AMUX = CLBLM_R_X15Y108_SLICE_X21Y108_AO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_DMUX = CLBLM_R_X15Y108_SLICE_X21Y108_DO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A = CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C = CLBLM_R_X15Y109_SLICE_X20Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D = CLBLM_R_X15Y109_SLICE_X20Y109_DO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_CMUX = CLBLM_R_X15Y109_SLICE_X20Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A = CLBLM_R_X15Y109_SLICE_X21Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B = CLBLM_R_X15Y109_SLICE_X21Y109_BO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C = CLBLM_R_X15Y109_SLICE_X21Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D = CLBLM_R_X15Y109_SLICE_X21Y109_DO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_AMUX = CLBLM_R_X15Y109_SLICE_X21Y109_AO5;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A = CLBLM_R_X15Y110_SLICE_X20Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C = CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D = CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_AMUX = CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A = CLBLM_R_X15Y110_SLICE_X21Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_AMUX = CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_BMUX = CLBLM_R_X15Y110_SLICE_X21Y110_BO5;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_CMUX = CLBLM_R_X15Y110_SLICE_X21Y110_CO5;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A = CLBLM_R_X15Y111_SLICE_X20Y111_AO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C = CLBLM_R_X15Y111_SLICE_X20Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D = CLBLM_R_X15Y111_SLICE_X20Y111_DO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_AMUX = CLBLM_R_X15Y111_SLICE_X20Y111_AO5;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_DMUX = CLBLM_R_X15Y111_SLICE_X20Y111_DO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A = CLBLM_R_X15Y111_SLICE_X21Y111_AO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B = CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C = CLBLM_R_X15Y111_SLICE_X21Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D = CLBLM_R_X15Y111_SLICE_X21Y111_DO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A = CLBLM_R_X15Y112_SLICE_X20Y112_AO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B = CLBLM_R_X15Y112_SLICE_X20Y112_BO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C = CLBLM_R_X15Y112_SLICE_X20Y112_CO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D = CLBLM_R_X15Y112_SLICE_X20Y112_DO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_AMUX = CLBLM_R_X15Y112_SLICE_X20Y112_AO5;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A = CLBLM_R_X15Y112_SLICE_X21Y112_AO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B = CLBLM_R_X15Y112_SLICE_X21Y112_BO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C = CLBLM_R_X15Y112_SLICE_X21Y112_CO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D = CLBLM_R_X15Y112_SLICE_X21Y112_DO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_BMUX = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_CMUX = CLBLM_R_X15Y112_SLICE_X21Y112_CO5;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A = CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B = CLBLM_R_X15Y113_SLICE_X20Y113_BO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C = CLBLM_R_X15Y113_SLICE_X20Y113_CO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D = CLBLM_R_X15Y113_SLICE_X20Y113_DO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C = CLBLM_R_X15Y113_SLICE_X21Y113_CO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D = CLBLM_R_X15Y113_SLICE_X21Y113_DO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A = CLBLM_R_X15Y114_SLICE_X20Y114_AO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B = CLBLM_R_X15Y114_SLICE_X20Y114_BO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C = CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_BMUX = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A = CLBLM_R_X15Y114_SLICE_X21Y114_AO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B = CLBLM_R_X15Y114_SLICE_X21Y114_BO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D = CLBLM_R_X15Y114_SLICE_X21Y114_DO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_BMUX = CLBLM_R_X15Y114_SLICE_X21Y114_BO5;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A = CLBLM_R_X15Y115_SLICE_X20Y115_AO6;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B = CLBLM_R_X15Y115_SLICE_X20Y115_BO6;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C = CLBLM_R_X15Y115_SLICE_X20Y115_CO6;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D = CLBLM_R_X15Y115_SLICE_X20Y115_DO6;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_BMUX = CLBLM_R_X15Y115_SLICE_X20Y115_BO5;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A = CLBLM_R_X15Y115_SLICE_X21Y115_AO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B = CLBLM_R_X15Y115_SLICE_X21Y115_BO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C = CLBLM_R_X15Y115_SLICE_X21Y115_CO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D = CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_CMUX = CLBLM_R_X15Y115_SLICE_X21Y115_CO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A = CLBLM_R_X15Y116_SLICE_X20Y116_AO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B = CLBLM_R_X15Y116_SLICE_X20Y116_BO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C = CLBLM_R_X15Y116_SLICE_X20Y116_CO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D = CLBLM_R_X15Y116_SLICE_X20Y116_DO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_CMUX = CLBLM_R_X15Y116_SLICE_X20Y116_CO5;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A = CLBLM_R_X15Y116_SLICE_X21Y116_AO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B = CLBLM_R_X15Y116_SLICE_X21Y116_BO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C = CLBLM_R_X15Y116_SLICE_X21Y116_CO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D = CLBLM_R_X15Y116_SLICE_X21Y116_DO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A = CLBLM_R_X15Y117_SLICE_X20Y117_AO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B = CLBLM_R_X15Y117_SLICE_X20Y117_BO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C = CLBLM_R_X15Y117_SLICE_X20Y117_CO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D = CLBLM_R_X15Y117_SLICE_X20Y117_DO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_BMUX = CLBLM_R_X15Y117_SLICE_X20Y117_BO5;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_CMUX = CLBLM_R_X15Y117_SLICE_X20Y117_CO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A = CLBLM_R_X15Y117_SLICE_X21Y117_AO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B = CLBLM_R_X15Y117_SLICE_X21Y117_BO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C = CLBLM_R_X15Y117_SLICE_X21Y117_CO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D = CLBLM_R_X15Y117_SLICE_X21Y117_DO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A = CLBLM_R_X15Y118_SLICE_X20Y118_AO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B = CLBLM_R_X15Y118_SLICE_X20Y118_BO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C = CLBLM_R_X15Y118_SLICE_X20Y118_CO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D = CLBLM_R_X15Y118_SLICE_X20Y118_DO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_BMUX = CLBLM_R_X15Y118_SLICE_X20Y118_BO5;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A = CLBLM_R_X15Y118_SLICE_X21Y118_AO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B = CLBLM_R_X15Y118_SLICE_X21Y118_BO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C = CLBLM_R_X15Y118_SLICE_X21Y118_CO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D = CLBLM_R_X15Y118_SLICE_X21Y118_DO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A = CLBLM_R_X15Y119_SLICE_X20Y119_AO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B = CLBLM_R_X15Y119_SLICE_X20Y119_BO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C = CLBLM_R_X15Y119_SLICE_X20Y119_CO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D = CLBLM_R_X15Y119_SLICE_X20Y119_DO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_BMUX = CLBLM_R_X15Y119_SLICE_X20Y119_BO5;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_CMUX = CLBLM_R_X15Y119_SLICE_X20Y119_CO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A = CLBLM_R_X15Y119_SLICE_X21Y119_AO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B = CLBLM_R_X15Y119_SLICE_X21Y119_BO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C = CLBLM_R_X15Y119_SLICE_X21Y119_CO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D = CLBLM_R_X15Y119_SLICE_X21Y119_DO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_CMUX = CLBLM_R_X15Y119_SLICE_X21Y119_CO5;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A = CLBLM_R_X15Y120_SLICE_X20Y120_AO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B = CLBLM_R_X15Y120_SLICE_X20Y120_BO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C = CLBLM_R_X15Y120_SLICE_X20Y120_CO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D = CLBLM_R_X15Y120_SLICE_X20Y120_DO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A = CLBLM_R_X15Y120_SLICE_X21Y120_AO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C = CLBLM_R_X15Y120_SLICE_X21Y120_CO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D = CLBLM_R_X15Y120_SLICE_X21Y120_DO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_BMUX = CLBLM_R_X15Y120_SLICE_X21Y120_BO5;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A = CLBLM_R_X15Y121_SLICE_X20Y121_AO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B = CLBLM_R_X15Y121_SLICE_X20Y121_BO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C = CLBLM_R_X15Y121_SLICE_X20Y121_CO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D = CLBLM_R_X15Y121_SLICE_X20Y121_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A = CLBLM_R_X15Y121_SLICE_X21Y121_AO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B = CLBLM_R_X15Y121_SLICE_X21Y121_BO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C = CLBLM_R_X15Y121_SLICE_X21Y121_CO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D = CLBLM_R_X15Y121_SLICE_X21Y121_DO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A = CLBLM_R_X15Y122_SLICE_X20Y122_AO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B = CLBLM_R_X15Y122_SLICE_X20Y122_BO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C = CLBLM_R_X15Y122_SLICE_X20Y122_CO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D = CLBLM_R_X15Y122_SLICE_X20Y122_DO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_CMUX = CLBLM_R_X15Y122_SLICE_X20Y122_CO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_DMUX = CLBLM_R_X15Y122_SLICE_X20Y122_DO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A = CLBLM_R_X15Y122_SLICE_X21Y122_AO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B = CLBLM_R_X15Y122_SLICE_X21Y122_BO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C = CLBLM_R_X15Y122_SLICE_X21Y122_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D = CLBLM_R_X15Y122_SLICE_X21Y122_DO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A = CLBLM_R_X15Y123_SLICE_X20Y123_AO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B = CLBLM_R_X15Y123_SLICE_X20Y123_BO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C = CLBLM_R_X15Y123_SLICE_X20Y123_CO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D = CLBLM_R_X15Y123_SLICE_X20Y123_DO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_BMUX = CLBLM_R_X15Y123_SLICE_X20Y123_BO5;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_CMUX = CLBLM_R_X15Y123_SLICE_X20Y123_CO5;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A = CLBLM_R_X15Y123_SLICE_X21Y123_AO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B = CLBLM_R_X15Y123_SLICE_X21Y123_BO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C = CLBLM_R_X15Y123_SLICE_X21Y123_CO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D = CLBLM_R_X15Y123_SLICE_X21Y123_DO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_BMUX = CLBLM_R_X15Y123_SLICE_X21Y123_BO5;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_CMUX = CLBLM_R_X15Y123_SLICE_X21Y123_CO5;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A = CLBLM_R_X15Y124_SLICE_X20Y124_AO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B = CLBLM_R_X15Y124_SLICE_X20Y124_BO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C = CLBLM_R_X15Y124_SLICE_X20Y124_CO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D = CLBLM_R_X15Y124_SLICE_X20Y124_DO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_BMUX = CLBLM_R_X15Y124_SLICE_X20Y124_BO5;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_CMUX = CLBLM_R_X15Y124_SLICE_X20Y124_CO5;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A = CLBLM_R_X15Y124_SLICE_X21Y124_AO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B = CLBLM_R_X15Y124_SLICE_X21Y124_BO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C = CLBLM_R_X15Y124_SLICE_X21Y124_CO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D = CLBLM_R_X15Y124_SLICE_X21Y124_DO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A = CLBLM_R_X15Y125_SLICE_X20Y125_AO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B = CLBLM_R_X15Y125_SLICE_X20Y125_BO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C = CLBLM_R_X15Y125_SLICE_X20Y125_CO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D = CLBLM_R_X15Y125_SLICE_X20Y125_DO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A = CLBLM_R_X15Y125_SLICE_X21Y125_AO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B = CLBLM_R_X15Y125_SLICE_X21Y125_BO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C = CLBLM_R_X15Y125_SLICE_X21Y125_CO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D = CLBLM_R_X15Y125_SLICE_X21Y125_DO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_CMUX = CLBLM_R_X15Y125_SLICE_X21Y125_CO5;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A = CLBLM_R_X15Y126_SLICE_X20Y126_AO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B = CLBLM_R_X15Y126_SLICE_X20Y126_BO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C = CLBLM_R_X15Y126_SLICE_X20Y126_CO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D = CLBLM_R_X15Y126_SLICE_X20Y126_DO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A = CLBLM_R_X15Y126_SLICE_X21Y126_AO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B = CLBLM_R_X15Y126_SLICE_X21Y126_BO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C = CLBLM_R_X15Y126_SLICE_X21Y126_CO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_DMUX = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A = CLBLM_R_X15Y127_SLICE_X20Y127_AO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B = CLBLM_R_X15Y127_SLICE_X20Y127_BO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C = CLBLM_R_X15Y127_SLICE_X20Y127_CO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D = CLBLM_R_X15Y127_SLICE_X20Y127_DO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A = CLBLM_R_X15Y127_SLICE_X21Y127_AO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_AMUX = CLBLM_R_X15Y127_SLICE_X21Y127_AO5;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B = CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_AMUX = CLBLM_R_X15Y128_SLICE_X20Y128_AO5;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_BMUX = CLBLM_R_X15Y128_SLICE_X20Y128_BO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A = CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D = CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_AMUX = CLBLM_R_X15Y128_SLICE_X21Y128_AO5;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A = CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B = CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C = CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D = CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A = CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C = CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_AMUX = CLBLM_R_X15Y129_SLICE_X21Y129_AO5;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_CMUX = CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A = CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B = CLBLM_R_X15Y130_SLICE_X20Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C = CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D = CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A = CLBLM_R_X15Y130_SLICE_X21Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B = CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C = CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D = CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A = CLBLM_R_X15Y131_SLICE_X20Y131_AO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B = CLBLM_R_X15Y131_SLICE_X20Y131_BO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C = CLBLM_R_X15Y131_SLICE_X20Y131_CO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D = CLBLM_R_X15Y131_SLICE_X20Y131_DO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_AMUX = CLBLM_R_X15Y131_SLICE_X20Y131_AO5;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_BMUX = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_CMUX = CLBLM_R_X15Y131_SLICE_X20Y131_CO5;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_DMUX = CLBLM_R_X15Y131_SLICE_X20Y131_DO5;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A = CLBLM_R_X15Y131_SLICE_X21Y131_AO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C = CLBLM_R_X15Y131_SLICE_X21Y131_CO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D = CLBLM_R_X15Y131_SLICE_X21Y131_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_AMUX = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A = CLBLM_R_X15Y132_SLICE_X20Y132_AO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B = CLBLM_R_X15Y132_SLICE_X20Y132_BO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C = CLBLM_R_X15Y132_SLICE_X20Y132_CO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D = CLBLM_R_X15Y132_SLICE_X20Y132_DO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A = CLBLM_R_X15Y132_SLICE_X21Y132_AO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B = CLBLM_R_X15Y132_SLICE_X21Y132_BO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C = CLBLM_R_X15Y132_SLICE_X21Y132_CO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D = CLBLM_R_X15Y132_SLICE_X21Y132_DO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_O = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_O = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_O = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_O = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_O = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_O = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_O = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_O = LIOB33_X0Y167_IOB_X0Y167_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_O = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_O = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_O = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_O = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_O = LIOB33_X0Y179_IOB_X0Y179_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_O = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_O = LIOB33_X0Y183_IOB_X0Y183_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_O = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_O = LIOB33_X0Y185_IOB_X0Y185_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_O = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_O = LIOB33_X0Y189_IOB_X0Y189_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_O = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_O = LIOB33_X0Y191_IOB_X0Y191_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_O = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_O = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_O = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_O = LIOB33_X0Y197_IOB_X0Y197_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_O = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_O = LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y144_D;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O = LIOB33_X0Y143_IOB_X0Y143_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O = LIOB33_X0Y169_IOB_X0Y169_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O = LIOB33_X0Y181_IOB_X0Y181_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O = LIOB33_X0Y193_IOB_X0Y193_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O = LIOB33_X0Y163_IOB_X0Y163_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O = LIOB33_X0Y187_IOB_X0Y187_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_OQ = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_OQ = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_OQ = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_OQ = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_OQ = CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_OQ = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = CLBLM_L_X16Y114_SLICE_X22Y114_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = CLBLM_R_X15Y114_SLICE_X21Y114_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLM_L_X16Y116_SLICE_X23Y116_AQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = CLBLM_L_X16Y114_SLICE_X23Y114_BQ;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLM_R_X15Y115_SLICE_X20Y115_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLM_R_X15Y116_SLICE_X20Y116_BQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLM_L_X16Y115_SLICE_X22Y115_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLM_R_X15Y115_SLICE_X21Y115_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLM_L_X16Y115_SLICE_X23Y115_BQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_L_X16Y115_SLICE_X23Y115_AQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_L_X16Y114_SLICE_X23Y114_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_R_X15Y116_SLICE_X21Y116_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_R_X15Y114_SLICE_X20Y114_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_R_X15Y117_SLICE_X21Y117_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_L_X16Y117_SLICE_X22Y117_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLM_R_X15Y119_SLICE_X20Y119_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLM_R_X15Y118_SLICE_X20Y118_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_L_X16Y119_SLICE_X22Y119_AQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_L_X16Y119_SLICE_X23Y119_AQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLM_R_X15Y132_SLICE_X21Y132_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLM_R_X15Y118_SLICE_X21Y118_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_R_X15Y132_SLICE_X21Y132_CQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLM_R_X15Y132_SLICE_X21Y132_BQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLM_R_X15Y132_SLICE_X21Y132_DQ;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_R_X15Y116_SLICE_X20Y116_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLM_L_X16Y116_SLICE_X23Y116_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_L_X16Y117_SLICE_X22Y117_AQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_R_X15Y116_SLICE_X21Y116_BQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLM_R_X15Y119_SLICE_X21Y119_BQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_R_X15Y119_SLICE_X21Y119_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_R_X15Y117_SLICE_X20Y117_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_R_X15Y117_SLICE_X21Y117_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLM_R_X15Y132_SLICE_X21Y132_DQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A3 = CLBLM_R_X15Y117_SLICE_X20Y117_CO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A4 = CLBLM_L_X16Y117_SLICE_X23Y117_AO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A5 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_A6 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B1 = CLBLM_R_X15Y117_SLICE_X21Y117_DO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B2 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B3 = CLBLM_L_X16Y116_SLICE_X22Y116_AO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B5 = CLBLM_L_X16Y117_SLICE_X22Y117_BQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_B6 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C1 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C2 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C3 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C4 = CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C5 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_C6 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D1 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D2 = CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D4 = CLBLM_R_X15Y117_SLICE_X21Y117_BQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_D6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y117_SLICE_X21Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A1 = CLBLM_R_X15Y117_SLICE_X20Y117_DO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A2 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A3 = CLBLM_R_X15Y118_SLICE_X20Y118_BO5;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A5 = CLBLM_R_X15Y117_SLICE_X21Y117_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B2 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B3 = CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B4 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B5 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_B6 = 1'b1;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C1 = CLBLM_R_X15Y117_SLICE_X21Y117_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C5 = CLBLM_R_X15Y117_SLICE_X20Y117_BO5;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_C6 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLM_R_X15Y119_SLICE_X20Y119_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D1 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D2 = CLBLM_R_X15Y117_SLICE_X20Y117_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_D6 = CLBLM_R_X15Y117_SLICE_X20Y117_BO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X15Y117_SLICE_X20Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y109_IOB_X1Y110_O = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLM_R_X15Y118_SLICE_X20Y118_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A2 = CLBLM_L_X12Y113_SLICE_X16Y113_BO5;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A3 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A4 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D4 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A1 = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A3 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A5 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B1 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B2 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B4 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B5 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B6 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C1 = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C2 = CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C3 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C6 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D1 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D2 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D4 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A1 = CLBLM_R_X15Y118_SLICE_X21Y118_DO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A3 = CLBLM_R_X15Y118_SLICE_X21Y118_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A4 = CLBLM_R_X15Y118_SLICE_X21Y118_BO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A5 = CLBLM_L_X16Y116_SLICE_X23Y116_DO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_A6 = CLBLM_R_X15Y119_SLICE_X21Y119_BQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B1 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B5 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_B6 = CLBLM_R_X15Y119_SLICE_X21Y119_CO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C1 = CLBLM_L_X16Y118_SLICE_X22Y118_AO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C4 = CLBLM_R_X15Y119_SLICE_X21Y119_BQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C5 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_C6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D1 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D5 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_D6 = CLBLM_L_X16Y118_SLICE_X22Y118_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y118_SLICE_X21Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A1 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A3 = CLBLM_R_X15Y117_SLICE_X20Y117_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A4 = CLBLM_R_X15Y118_SLICE_X20Y118_BO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_A6 = CLBLM_R_X15Y118_SLICE_X20Y118_CO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B2 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B3 = CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B4 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B5 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_B6 = 1'b1;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C2 = CLBLM_R_X15Y118_SLICE_X20Y118_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C4 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C5 = CLBLM_R_X15Y118_SLICE_X20Y118_DO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_C6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D1 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D2 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D3 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D4 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D5 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_D6 = CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  assign CLBLM_R_X15Y118_SLICE_X20Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A1 = CLBLM_L_X12Y115_SLICE_X16Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A3 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A4 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A6 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_AX = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B2 = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B3 = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B4 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B5 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C1 = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C4 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C5 = CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A1 = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A3 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A4 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A5 = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B1 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B2 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B3 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B4 = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B5 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C3 = CLBLM_L_X12Y115_SLICE_X16Y115_A5Q;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C4 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C5 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C6 = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D3 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D4 = CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D5 = CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A1 = CLBLM_R_X15Y119_SLICE_X21Y119_DO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A2 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A3 = CLBLM_L_X16Y119_SLICE_X22Y119_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A5 = CLBLM_R_X15Y119_SLICE_X21Y119_CO5;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_A6 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B1 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B3 = CLBLM_R_X15Y119_SLICE_X21Y119_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B4 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B5 = CLBLM_R_X15Y118_SLICE_X21Y118_CO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_B6 = CLBLM_R_X15Y119_SLICE_X21Y119_CO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C1 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C2 = CLBLM_R_X15Y117_SLICE_X21Y117_CO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C3 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C4 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C5 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_C6 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D2 = CLBLM_R_X15Y119_SLICE_X21Y119_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D3 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D5 = CLBLM_L_X16Y119_SLICE_X22Y119_CO6;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_D6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y119_SLICE_X21Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A1 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A3 = CLBLM_R_X15Y118_SLICE_X20Y118_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A5 = CLBLM_R_X15Y119_SLICE_X20Y119_CO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_A6 = CLBLM_R_X15Y117_SLICE_X21Y117_CO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B1 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B2 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B3 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B4 = CLBLM_R_X15Y118_SLICE_X20Y118_DO6;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B5 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_B6 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C2 = CLBLM_R_X15Y119_SLICE_X20Y119_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C3 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C5 = CLBLM_R_X15Y119_SLICE_X20Y119_BO5;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_C6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D1 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D2 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D3 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D4 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D5 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_D6 = 1'b1;
  assign CLBLM_R_X15Y119_SLICE_X20Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A2 = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A3 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A5 = CLBLM_L_X12Y116_SLICE_X17Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_A6 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_L_X16Y119_SLICE_X22Y119_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B1 = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B3 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_B6 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C1 = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C3 = CLBLM_L_X12Y116_SLICE_X16Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C4 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_L_X16Y119_SLICE_X23Y119_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D1 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D2 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D3 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D4 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D5 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_D6 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X17Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A1 = CLBLM_L_X12Y116_SLICE_X16Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A5 = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_A6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B1 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B2 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_B6 = 1'b1;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C1 = CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C3 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C4 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_C6 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D2 = CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D3 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D4 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D5 = CLBLM_L_X12Y116_SLICE_X16Y116_BO5;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y116_SLICE_X16Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A1 = CLBLM_R_X15Y120_SLICE_X21Y120_BO5;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A2 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A3 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A4 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_A6 = CLBLM_R_X15Y121_SLICE_X21Y121_CO6;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_B6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C1 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C2 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C3 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C4 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C5 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_C6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D1 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D2 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D3 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D4 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A1 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A2 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A3 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A4 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_A6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_D6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A1 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B1 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B2 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B3 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B4 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_B6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A2 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A4 = CLBLM_R_X15Y120_SLICE_X20Y120_BO6;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C1 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C2 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C3 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C4 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_C6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B1 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B3 = CLBLM_R_X15Y120_SLICE_X20Y120_AQ;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B5 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_B6 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D1 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D2 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D3 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B5 = CLBLM_L_X16Y107_SLICE_X23Y107_DO5;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D4 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X15Y100_D6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B6 = CLBLM_L_X16Y108_SLICE_X22Y108_CO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A2 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_A6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D2 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D3 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D4 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B2 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B5 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_B6 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C1 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C2 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C4 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C5 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_C6 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D1 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D2 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D3 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D4 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D5 = 1'b1;
  assign CLBLM_R_X11Y100_SLICE_X14Y100_D6 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A2 = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A4 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A5 = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A6 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B1 = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B2 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B3 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B4 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B5 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C1 = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C4 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C5 = CLBLM_L_X12Y116_SLICE_X17Y116_BO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D4 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A1 = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A2 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A4 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B1 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B2 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B5 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C2 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C4 = CLBLM_L_X12Y116_SLICE_X17Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C5 = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C6 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D2 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D4 = CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D5 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A1 = CLBLM_R_X15Y121_SLICE_X21Y121_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A4 = CLBLM_L_X16Y121_SLICE_X22Y121_AQ;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A5 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_A6 = CLBLM_R_X15Y124_SLICE_X20Y124_CO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B1 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B3 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B5 = CLBLM_L_X16Y121_SLICE_X22Y121_AQ;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C1 = CLBLM_R_X15Y120_SLICE_X21Y120_AQ;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C2 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C5 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_C6 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D1 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D3 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D5 = CLBLM_R_X15Y121_SLICE_X21Y121_AQ;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A1 = 1'b1;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A3 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A4 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A5 = 1'b1;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_A6 = 1'b1;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_D6 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A1 = CLBLM_R_X15Y121_SLICE_X20Y121_DO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B1 = CLBLM_R_X11Y100_SLICE_X14Y100_CO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B2 = CLBLM_R_X11Y102_SLICE_X14Y102_AO5;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B3 = CLBLM_R_X11Y100_SLICE_X14Y100_AO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B4 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B5 = CLBLM_R_X11Y101_SLICE_X15Y101_AO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_B6 = CLBLM_R_X11Y101_SLICE_X15Y101_AO5;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A2 = CLBLM_R_X15Y123_SLICE_X20Y123_AQ;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C1 = CLBLM_R_X11Y101_SLICE_X15Y101_AO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C3 = CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_C6 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B1 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B4 = CLBLM_R_X15Y120_SLICE_X20Y120_AQ;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B5 = CLBLM_R_X15Y124_SLICE_X20Y124_BO5;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_B6 = CLBLM_R_X15Y121_SLICE_X20Y121_CO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D1 = 1'b1;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D2 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D3 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D4 = CLBLM_R_X11Y102_SLICE_X14Y102_AO5;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D5 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y101_SLICE_X15Y101_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C6 = CLBLM_R_X15Y121_SLICE_X20Y121_BQ;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A1 = 1'b1;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A2 = CLBLM_R_X11Y101_SLICE_X15Y101_DO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A3 = CLBLM_R_X11Y103_SLICE_X14Y103_CO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A5 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_A6 = CLBLM_R_X11Y101_SLICE_X14Y101_CO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D2 = CLBLM_R_X15Y121_SLICE_X20Y121_AQ;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D3 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D4 = CLBLM_R_X15Y120_SLICE_X20Y120_CO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D5 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B1 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B2 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B3 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_B6 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C2 = CLBLM_R_X11Y102_SLICE_X14Y102_AO5;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C3 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C4 = CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C5 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_C6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D1 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D2 = CLBLM_R_X11Y100_SLICE_X14Y100_AO5;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D3 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D4 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D5 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_D6 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X11Y101_SLICE_X14Y101_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLM_R_X15Y132_SLICE_X21Y132_AQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A2 = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A4 = CLBLM_R_X15Y122_SLICE_X21Y122_BO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A5 = CLBLM_R_X15Y123_SLICE_X21Y123_AQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B1 = CLBLM_R_X15Y122_SLICE_X21Y122_DO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B2 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B3 = CLBLM_R_X15Y122_SLICE_X21Y122_AQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_B6 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLM_R_X15Y118_SLICE_X21Y118_AQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C1 = CLBLM_R_X15Y122_SLICE_X20Y122_AQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C2 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C5 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A1 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A2 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A3 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_A6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A1 = CLBLM_R_X15Y122_SLICE_X21Y122_CO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B1 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B2 = CLBLM_L_X12Y102_SLICE_X17Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B3 = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B4 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B5 = CLBLM_R_X11Y102_SLICE_X15Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_B6 = CLBLM_R_X11Y102_SLICE_X15Y102_AO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A2 = CLBLM_R_X15Y122_SLICE_X20Y122_BQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A3 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B1 = CLBLM_R_X15Y123_SLICE_X20Y123_BO5;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C1 = CLBLM_R_X11Y102_SLICE_X15Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C4 = CLBLM_R_X11Y103_SLICE_X15Y103_BO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C5 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_C6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B3 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B4 = CLBLM_R_X15Y122_SLICE_X20Y122_DO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B5 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_B6 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D1 = CLBLM_L_X12Y102_SLICE_X17Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D2 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D3 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D4 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D5 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X15Y102_D6 = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D1 = CLBLM_R_X15Y122_SLICE_X20Y122_BQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A2 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A3 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A5 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_A6 = 1'b1;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D2 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D3 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D4 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B1 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B2 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B3 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B4 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_B6 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C1 = CLBLM_L_X12Y102_SLICE_X17Y102_AO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C2 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C4 = CLBLM_R_X11Y100_SLICE_X14Y100_CO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C5 = CLBLM_R_X11Y102_SLICE_X14Y102_DO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_C6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D1 = CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D2 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D3 = 1'b1;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y102_SLICE_X14Y102_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A1 = CLBLM_R_X15Y123_SLICE_X21Y123_DO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A2 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A3 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A5 = CLBLM_R_X15Y123_SLICE_X21Y123_CO5;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_A6 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_B6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_C6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D1 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D2 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D3 = CLBLM_R_X15Y123_SLICE_X21Y123_AQ;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A1 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A2 = CLBLM_R_X11Y102_SLICE_X15Y102_DO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A3 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_D6 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A1 = CLBLM_R_X15Y123_SLICE_X20Y123_DO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B1 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B2 = CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B3 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B4 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B5 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B6 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A2 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A3 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A4 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C1 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C2 = CLBLM_R_X11Y102_SLICE_X15Y102_DO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_B6 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D1 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D3 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D5 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A1 = CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A3 = CLBLM_R_X11Y103_SLICE_X15Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A4 = CLBLM_R_X11Y103_SLICE_X14Y103_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A5 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D3 = CLBLM_R_X15Y123_SLICE_X20Y123_AQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D4 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B1 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B2 = CLBLM_R_X11Y102_SLICE_X14Y102_AO5;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B3 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B5 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C2 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C3 = CLBLM_R_X11Y103_SLICE_X15Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C6 = CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D1 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D3 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A1 = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A2 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A4 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B1 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C4 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C5 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D2 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A1 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A2 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A4 = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A6 = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C1 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C2 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C4 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D2 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D3 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D4 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A1 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A3 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A4 = CLBLM_R_X15Y124_SLICE_X21Y124_BO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_A6 = CLBLM_R_X15Y123_SLICE_X21Y123_CO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B1 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B2 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B3 = CLBLM_R_X15Y124_SLICE_X21Y124_AQ;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_B6 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C1 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C4 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C5 = CLBLM_R_X15Y125_SLICE_X21Y125_BQ;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D2 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D3 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D4 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A3 = CLBLM_R_X11Y103_SLICE_X15Y103_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A5 = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A6 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_D6 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A1 = CLBLM_R_X15Y124_SLICE_X20Y124_DO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B6 = 1'b1;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A4 = CLBLM_R_X15Y127_SLICE_X20Y127_AQ;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C6 = 1'b1;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C3 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D6 = 1'b1;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_C6 = 1'b1;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A1 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A2 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A4 = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A6 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D5 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_D6 = CLBLM_R_X15Y124_SLICE_X20Y124_AQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B1 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B3 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_R_X15Y132_SLICE_X21Y132_CQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C3 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C4 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C5 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D1 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D3 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D6 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLM_R_X15Y132_SLICE_X21Y132_BQ;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A1 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A4 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B3 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C2 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C3 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D6 = 1'b1;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A1 = CLBLM_R_X15Y125_SLICE_X21Y125_DO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A2 = CLBLM_R_X15Y126_SLICE_X21Y126_AQ;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A3 = CLBLM_R_X15Y123_SLICE_X21Y123_BO5;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B1 = CLBLM_R_X15Y125_SLICE_X21Y125_AQ;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B4 = CLBLM_R_X15Y124_SLICE_X21Y124_CO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B5 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_B6 = CLBLM_R_X15Y125_SLICE_X21Y125_CO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_C6 = 1'b1;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D1 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D4 = CLBLM_R_X15Y125_SLICE_X21Y125_AQ;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D5 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_D6 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A1 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A3 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A4 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A5 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B2 = CLBLM_R_X15Y124_SLICE_X21Y124_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B3 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B4 = CLBLM_R_X15Y126_SLICE_X20Y126_BQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B5 = CLBLM_R_X15Y130_SLICE_X20Y130_BQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_B6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C1 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C2 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C4 = 1'b1;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C5 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D1 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D2 = CLBLM_R_X15Y126_SLICE_X20Y126_BQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D4 = 1'b1;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D5 = CLBLM_R_X15Y124_SLICE_X21Y124_AQ;
  assign CLBLM_R_X15Y125_SLICE_X20Y125_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B6 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C4 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C5 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A1 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A4 = CLBLM_L_X12Y122_SLICE_X17Y122_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B2 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_B6 = CLBLM_L_X12Y122_SLICE_X17Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C2 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C3 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C4 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_C6 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D4 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D2 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A1 = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A3 = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A4 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A5 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A6 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y122_SLICE_X17Y122_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A1 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B1 = CLBLM_L_X10Y101_SLICE_X13Y101_AO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B3 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B4 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A4 = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A5 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A6 = CLBLM_L_X12Y122_SLICE_X16Y122_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C1 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C3 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B2 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B3 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C6 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B4 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B5 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D2 = CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D4 = CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D5 = 1'b1;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D1 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D2 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A2 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A3 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A4 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A5 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A6 = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D3 = CLBLM_L_X12Y121_SLICE_X17Y121_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D5 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B1 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B2 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B3 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B5 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B6 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C1 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C4 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C5 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C6 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D1 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D2 = CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D3 = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D4 = CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D5 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D6 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A1 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A3 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A4 = CLBLM_R_X15Y126_SLICE_X21Y126_BO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A5 = CLBLM_R_X15Y124_SLICE_X21Y124_AQ;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_A6 = CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B1 = CLBLM_R_X15Y126_SLICE_X21Y126_AQ;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B2 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B3 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C1 = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C3 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C5 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_C6 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D4 = CLBLM_R_X15Y126_SLICE_X21Y126_CO6;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D5 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_D6 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A1 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A2 = CLBLM_R_X15Y126_SLICE_X20Y126_BQ;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A3 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B1 = CLBLM_R_X15Y126_SLICE_X20Y126_DO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B3 = CLBLM_R_X15Y123_SLICE_X20Y123_CO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B4 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_B6 = CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C4 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D1 = CLBLM_R_X15Y126_SLICE_X20Y126_BQ;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D2 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_D6 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A1 = CLBLM_L_X12Y123_SLICE_X17Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A3 = CLBLM_L_X12Y122_SLICE_X17Y122_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A5 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B4 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B5 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_B6 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C4 = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_C6 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D1 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D2 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D3 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A2 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A4 = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A6 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D5 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_D6 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B1 = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B3 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B4 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A2 = CLBLM_L_X12Y123_SLICE_X17Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C4 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C5 = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C6 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B1 = CLBLM_L_X12Y123_SLICE_X16Y123_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B4 = CLBLM_R_X15Y121_SLICE_X21Y121_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B5 = CLBLM_L_X12Y123_SLICE_X16Y123_CO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D1 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D6 = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A2 = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A5 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A6 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D2 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D4 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D5 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B3 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B4 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B5 = CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B6 = 1'b1;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C1 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C2 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C5 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D4 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D5 = CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D6 = 1'b1;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_A6 = 1'b1;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B2 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B3 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B4 = CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C2 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C3 = CLBLM_R_X15Y127_SLICE_X20Y127_DO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D2 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D3 = CLBLM_R_X15Y128_SLICE_X21Y128_AO5;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D4 = CLBLM_R_X15Y127_SLICE_X21Y127_AO5;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D5 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = 1'b1;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_D6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = 1'b1;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A3 = CLBLM_R_X15Y126_SLICE_X20Y126_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A4 = CLBLM_R_X15Y127_SLICE_X20Y127_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = 1'b1;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B1 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B2 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B3 = CLBLM_R_X15Y127_SLICE_X20Y127_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B4 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B5 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_B6 = CLBLM_R_X15Y127_SLICE_X20Y127_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = 1'b1;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D2 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D3 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A1 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A2 = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A4 = CLBLM_L_X12Y124_SLICE_X17Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_A6 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B4 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_B6 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C3 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C4 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_C6 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D3 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D4 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D5 = CLBLM_L_X12Y123_SLICE_X16Y123_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_D6 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y124_SLICE_X17Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A2 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A3 = CLBLM_L_X12Y123_SLICE_X16Y123_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B1 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B2 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B3 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B5 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_B6 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C3 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C6 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = 1'b1;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D4 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B1 = CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B5 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C1 = CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C2 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C3 = CLBLM_R_X15Y128_SLICE_X20Y128_BO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C4 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C6 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D2 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D4 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D6 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A2 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C4 = CLBLM_R_X15Y128_SLICE_X20Y128_AO5;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D3 = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D4 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A2 = CLBLM_R_X15Y127_SLICE_X20Y127_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A4 = CLBLM_R_X15Y125_SLICE_X21Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_A6 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B1 = CLBLM_L_X12Y125_SLICE_X17Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B2 = CLBLM_R_X15Y127_SLICE_X20Y127_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_B6 = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C3 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C4 = CLBLM_R_X15Y125_SLICE_X20Y125_CO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_C6 = CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D1 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D4 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_L_X12Y125_SLICE_X17Y125_D6 = CLBLM_R_X15Y125_SLICE_X21Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A1 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A2 = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A4 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B1 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B3 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B4 = CLBLM_L_X12Y125_SLICE_X16Y125_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C3 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D1 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D2 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D3 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B4 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B6 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C4 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D1 = CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D2 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A2 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A3 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A4 = CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B2 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B3 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B4 = CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B5 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B6 = CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D5 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A2 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A4 = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A5 = CLBLM_R_X15Y124_SLICE_X20Y124_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A6 = CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B2 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B3 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B4 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B5 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B6 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D2 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D3 = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D4 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D6 = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A2 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C3 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D3 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D5 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A1 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A4 = CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A6 = CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B2 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C2 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C3 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C4 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C5 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D6 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A1 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B1 = CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B4 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C3 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C4 = CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C6 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D3 = CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D4 = CLBLM_R_X15Y130_SLICE_X20Y130_BQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A2 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A4 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A5 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A6 = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B2 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B5 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B6 = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D1 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D5 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D6 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A1 = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A2 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B1 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B2 = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B3 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B4 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B6 = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D2 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D4 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D5 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y115_IOB_X1Y116_O = CLBLM_L_X16Y114_SLICE_X22Y114_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A1 = CLBLM_R_X15Y131_SLICE_X20Y131_CO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A3 = CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A4 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A6 = CLBLM_R_X15Y132_SLICE_X21Y132_DQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_AX = CLBLM_R_X15Y131_SLICE_X20Y131_AO5;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B1 = CLBLM_R_X15Y131_SLICE_X20Y131_CO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_BQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B5 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B6 = CLBLM_R_X15Y131_SLICE_X20Y131_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C1 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C2 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C3 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C4 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C5 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D1 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D2 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D3 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D4 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A2 = CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A4 = CLBLM_R_X15Y131_SLICE_X20Y131_DO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B1 = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B5 = CLBLM_R_X15Y131_SLICE_X20Y131_CO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C3 = CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C4 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D2 = CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D4 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D5 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_T1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A2 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A4 = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A5 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A6 = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C2 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C3 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C4 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C6 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D2 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D4 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D6 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A1 = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A2 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A3 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B1 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B2 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B4 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D1 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D2 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D3 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A3 = CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A5 = CLBLM_R_X15Y118_SLICE_X21Y118_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_A6 = CLBLM_R_X15Y132_SLICE_X21Y132_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B2 = CLBLM_R_X15Y132_SLICE_X21Y132_BQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_BQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_B6 = CLBLM_R_X15Y132_SLICE_X21Y132_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C2 = CLBLM_R_X15Y132_SLICE_X21Y132_CQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C4 = CLBLM_R_X15Y132_SLICE_X21Y132_BQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C5 = CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D2 = CLBLM_R_X15Y132_SLICE_X21Y132_CQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D3 = CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D4 = CLBLM_R_X15Y132_SLICE_X21Y132_DQ;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A1 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A4 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A6 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_D6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B1 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B2 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B5 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B6 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C2 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C3 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C4 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B2 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B4 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D1 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D2 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D3 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D6 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D1 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A3 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A4 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A5 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A6 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D3 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D4 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B1 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B3 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B5 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B6 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C1 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C2 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C2 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C4 = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C5 = CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C6 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D4 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D5 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A1 = CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A2 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B3 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C4 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C6 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D1 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D3 = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A1 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A6 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B2 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B4 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B5 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B6 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A5 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B3 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B5 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B6 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = CLBLM_L_X12Y116_SLICE_X16Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C5 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C6 = CLBLM_R_X15Y126_SLICE_X20Y126_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A1 = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A3 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B5 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B6 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C2 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C3 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C4 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D2 = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D3 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A1 = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A5 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B3 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B5 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C2 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C3 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C5 = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C6 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D2 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D4 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D5 = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = CLBLM_L_X12Y125_SLICE_X17Y125_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_AX = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = CLBLM_R_X13Y124_SLICE_X18Y124_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_R_X13Y124_SLICE_X18Y124_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = CLBLM_L_X12Y125_SLICE_X17Y125_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = CLBLM_R_X13Y121_SLICE_X18Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = CLBLM_L_X12Y123_SLICE_X16Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = CLBLM_R_X15Y120_SLICE_X21Y120_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = CLBLM_L_X12Y124_SLICE_X16Y124_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = CLBLM_L_X12Y124_SLICE_X16Y124_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = CLBLM_R_X13Y121_SLICE_X18Y121_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = CLBLM_R_X13Y125_SLICE_X19Y125_BO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = CLBLM_L_X12Y124_SLICE_X17Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = CLBLM_L_X16Y126_SLICE_X22Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = CLBLM_L_X16Y126_SLICE_X22Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = CLBLM_R_X13Y125_SLICE_X19Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLM_R_X15Y132_SLICE_X21Y132_DQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A1 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A2 = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A4 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A5 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A6 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B2 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B4 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B5 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C1 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C2 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C3 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C6 = CLBLM_L_X12Y126_SLICE_X17Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D1 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D2 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D3 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D6 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A3 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B4 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C3 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C6 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A1 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A2 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A3 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A4 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A5 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_A6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B1 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B2 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B3 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B4 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B5 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_B6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C1 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C2 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C3 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C4 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C5 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_C6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D1 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D2 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D3 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D4 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D5 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X23Y101_D6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A1 = CLBLM_L_X16Y101_SLICE_X22Y101_DO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A3 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A4 = CLBLM_R_X15Y103_SLICE_X21Y103_BO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A5 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_A6 = CLBLM_L_X16Y101_SLICE_X22Y101_CO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B1 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B2 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B4 = CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B5 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_B6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C1 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C2 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C4 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C5 = CLBLM_L_X16Y101_SLICE_X22Y101_BO5;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_C6 = CLBLM_L_X16Y102_SLICE_X22Y102_BO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D1 = CLBLM_R_X15Y100_SLICE_X21Y100_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D5 = CLBLM_L_X16Y102_SLICE_X22Y102_CO6;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C1 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C3 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C4 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C6 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D1 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D3 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D6 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A1 = CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A4 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B1 = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B3 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B4 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B6 = CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C4 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D2 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D3 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D4 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D5 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D6 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A1 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A2 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A5 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_A6 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B1 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B2 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B3 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B4 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B5 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_B6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C1 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C2 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C3 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C4 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C5 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_C6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D1 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D2 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D3 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D4 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D5 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X23Y102_D6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A1 = CLBLM_L_X16Y102_SLICE_X22Y102_DO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A2 = CLBLM_L_X16Y103_SLICE_X22Y103_BO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A4 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A5 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_A6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B1 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B2 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B4 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B5 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_B6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C2 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C3 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C4 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C5 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_C6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = 1'b1;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D3 = CLBLM_R_X15Y103_SLICE_X21Y103_AO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D1 = CLBLM_L_X16Y101_SLICE_X22Y101_BO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D6 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D2 = CLBLM_L_X16Y102_SLICE_X23Y102_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A1 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A2 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A3 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A4 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A5 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_A6 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B1 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B4 = CLBLM_L_X16Y102_SLICE_X23Y102_AO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B5 = CLBLM_R_X15Y108_SLICE_X21Y108_AO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_B6 = CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C2 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C3 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C4 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C5 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_C6 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D1 = CLBLM_L_X16Y103_SLICE_X23Y103_AO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D2 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D3 = CLBLM_R_X15Y100_SLICE_X21Y100_AO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X16Y103_SLICE_X23Y103_D6 = 1'b1;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A1 = CLBLM_R_X15Y103_SLICE_X21Y103_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A2 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A4 = CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_A6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B2 = CLBLM_L_X16Y103_SLICE_X23Y103_BO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B3 = CLBLM_R_X15Y103_SLICE_X20Y103_AO5;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B4 = CLBLM_R_X15Y103_SLICE_X21Y103_DO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B5 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C1 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C2 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C3 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C4 = CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C5 = CLBLM_L_X16Y102_SLICE_X22Y102_CO5;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D1 = 1'b1;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D2 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D3 = CLBLM_R_X15Y103_SLICE_X21Y103_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D4 = 1'b1;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D5 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A1 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A3 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A5 = CLBLM_R_X15Y129_SLICE_X21Y129_AO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A6 = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B2 = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B3 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B4 = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B5 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B6 = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C1 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C4 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C5 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D1 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D3 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D4 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D5 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A1 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A3 = CLBLM_L_X12Y124_SLICE_X16Y124_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A4 = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C3 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D1 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D5 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D6 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y120_SLICE_X21Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A2 = 1'b1;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A3 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A4 = CLBLM_L_X16Y104_SLICE_X23Y104_BO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A5 = 1'b1;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_A6 = CLBLM_R_X15Y106_SLICE_X20Y106_CO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A5 = CLBLM_R_X15Y123_SLICE_X21Y123_BO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B1 = CLBLM_L_X16Y103_SLICE_X23Y103_DO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B3 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B5 = CLBLM_L_X16Y105_SLICE_X23Y105_AO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_B6 = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_A6 = CLBLM_R_X15Y121_SLICE_X20Y121_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C1 = CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C2 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C3 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C4 = CLBLM_L_X16Y102_SLICE_X22Y102_CO5;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C5 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_C6 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = 1'b0;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D1 = CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D2 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D3 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D4 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D5 = CLBLM_L_X16Y102_SLICE_X22Y102_CO5;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_D6 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y104_SLICE_X23Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A2 = CLBLM_L_X16Y104_SLICE_X22Y104_DO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A4 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A5 = CLBLM_L_X16Y103_SLICE_X22Y103_DO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_A6 = CLBLM_R_X15Y104_SLICE_X21Y104_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_D6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = CLBLM_L_X12Y125_SLICE_X16Y125_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C2 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C5 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A1 = CLBLM_R_X15Y100_SLICE_X21Y100_DO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A2 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A3 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A4 = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_A6 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B1 = CLBLM_R_X15Y100_SLICE_X21Y100_DO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B2 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B3 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B4 = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_B6 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C1 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C2 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C3 = CLBLM_L_X16Y102_SLICE_X22Y102_BO5;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C4 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C5 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_C6 = CLBLM_R_X15Y103_SLICE_X20Y103_DO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D1 = CLBLM_R_X15Y103_SLICE_X20Y103_DO6;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D2 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D3 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D4 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D5 = CLBLM_L_X16Y102_SLICE_X22Y102_BO5;
  assign CLBLM_L_X16Y105_SLICE_X23Y105_D6 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D2 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A1 = CLBLM_L_X16Y105_SLICE_X22Y105_DO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A2 = CLBLM_L_X16Y104_SLICE_X23Y104_CO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A3 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A4 = CLBLM_L_X16Y105_SLICE_X22Y105_BO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B1 = CLBLM_L_X16Y108_SLICE_X22Y108_AO5;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A1 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A2 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A3 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A4 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A5 = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B1 = CLBLM_R_X15Y100_SLICE_X21Y100_AO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B2 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B3 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B4 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B5 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_B6 = 1'b1;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C1 = CLBLM_L_X16Y106_SLICE_X23Y106_AO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C3 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C4 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_C6 = CLBLM_L_X16Y105_SLICE_X23Y105_BO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D1 = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D2 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D3 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D4 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y106_SLICE_X23Y106_D6 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A1 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A3 = CLBLM_L_X16Y106_SLICE_X23Y106_CO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A4 = 1'b1;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A5 = CLBLM_L_X16Y106_SLICE_X22Y106_CO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_A6 = CLBLM_R_X15Y106_SLICE_X21Y106_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B1 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B2 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = LIOB33_X0Y187_IOB_X0Y188_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B5 = CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C5 = CLBLM_L_X16Y106_SLICE_X22Y106_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D1 = CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D2 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D3 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A1 = CLBLM_L_X16Y106_SLICE_X23Y106_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A3 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A5 = CLBLM_L_X16Y107_SLICE_X23Y107_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_A6 = CLBLM_L_X16Y107_SLICE_X23Y107_CO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B2 = CLBLM_L_X16Y110_SLICE_X23Y110_BO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B3 = CLBLM_L_X16Y106_SLICE_X23Y106_BO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B4 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_B6 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C1 = CLBLM_L_X16Y106_SLICE_X22Y106_BO5;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C2 = CLBLM_L_X16Y106_SLICE_X23Y106_BO5;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C5 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_C6 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D1 = CLBLM_L_X16Y105_SLICE_X23Y105_BO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D2 = CLBLM_L_X16Y106_SLICE_X22Y106_BO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D3 = CLBLM_L_X16Y106_SLICE_X23Y106_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D4 = CLBLM_L_X16Y105_SLICE_X23Y105_DO6;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D5 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X23Y107_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A1 = CLBLM_L_X16Y107_SLICE_X22Y107_DO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A2 = CLBLM_L_X16Y107_SLICE_X23Y107_DO5;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A3 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A4 = CLBLM_L_X16Y107_SLICE_X22Y107_BO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B1 = CLBLM_L_X16Y104_SLICE_X23Y104_DO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B5 = CLBLM_L_X16Y108_SLICE_X23Y108_AO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B6 = CLBLM_L_X16Y106_SLICE_X23Y106_AO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C5 = CLBLM_L_X16Y104_SLICE_X23Y104_DO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D2 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D3 = CLBLM_R_X15Y107_SLICE_X21Y107_AO5;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D4 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D5 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B2 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B4 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C2 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C4 = CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C5 = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A1 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A2 = CLBLM_L_X16Y110_SLICE_X23Y110_BO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A3 = CLBLM_L_X16Y108_SLICE_X22Y108_AO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A4 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A5 = CLBLM_L_X16Y109_SLICE_X23Y109_AO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B1 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B2 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B3 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B4 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B5 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_B6 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D5 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C1 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C2 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C3 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C4 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C5 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_C6 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D1 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D2 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D3 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D4 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D5 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X23Y108_D6 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A2 = CLBLM_L_X16Y109_SLICE_X22Y109_BO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A3 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A4 = CLBLM_L_X16Y109_SLICE_X22Y109_AO5;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A5 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = 1'b1;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B3 = CLBLM_L_X16Y107_SLICE_X22Y107_CO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B4 = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C1 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C3 = CLBLM_R_X15Y107_SLICE_X21Y107_AO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_C6 = CLBLM_L_X16Y106_SLICE_X22Y106_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D1 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D5 = CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D6 = CLBLM_R_X15Y108_SLICE_X20Y108_AO6;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_D3 = CLBLM_R_X15Y108_SLICE_X21Y108_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y108_SLICE_X22Y108_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign CLBLM_R_X15Y121_SLICE_X21Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A1 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A2 = CLBLM_L_X16Y110_SLICE_X22Y110_BO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A3 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A4 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A5 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_A6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_B6 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A5 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C1 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C2 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C3 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C4 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C5 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_C6 = CLBLM_L_X16Y110_SLICE_X22Y110_BO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_A6 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_D1 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D1 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D2 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D3 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D4 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D5 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X23Y109_D6 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A1 = CLBLM_L_X16Y109_SLICE_X22Y109_BO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A2 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A3 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A4 = CLBLM_L_X16Y110_SLICE_X22Y110_BO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A5 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B1 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B2 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B3 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B4 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_B5 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = 1'b1;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C1 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C2 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C3 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_C6 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D1 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D2 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D3 = CLBLM_R_X15Y107_SLICE_X21Y107_CQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D5 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y109_SLICE_X22Y109_D6 = CLBLM_L_X16Y110_SLICE_X22Y110_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C1 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_C5 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A5 = CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A6 = CLBLM_R_X13Y123_SLICE_X18Y123_CO6;
  assign CLBLM_R_X15Y121_SLICE_X20Y121_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C1 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C2 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C5 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A3 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_A6 = 1'b1;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B3 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C2 = 1'b1;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C3 = CLBLM_L_X16Y109_SLICE_X23Y109_AO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C4 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_C6 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D3 = 1'b1;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D4 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X23Y110_D6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A1 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A2 = CLBLM_L_X16Y109_SLICE_X22Y109_CO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A4 = CLBLM_R_X15Y111_SLICE_X20Y111_DO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_A6 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B2 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B3 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B4 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B5 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_B6 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C1 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C4 = CLBLM_L_X16Y109_SLICE_X22Y109_AO5;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C5 = 1'b1;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D6 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D1 = 1'b1;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D3 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_D6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X16Y110_SLICE_X22Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A1 = CLBLM_R_X15Y111_SLICE_X20Y111_BO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A2 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A3 = CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A4 = CLBLM_L_X16Y111_SLICE_X23Y111_BO6;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A5 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B1 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_B6 = 1'b1;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C1 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C2 = CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C3 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C4 = CLBLM_R_X15Y110_SLICE_X21Y110_BO5;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C5 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_C6 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D1 = CLBLM_R_X15Y110_SLICE_X21Y110_BO5;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D2 = CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D3 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D4 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D5 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_D6 = 1'b1;
  assign CLBLM_L_X16Y111_SLICE_X23Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A1 = CLBLM_L_X16Y110_SLICE_X23Y110_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A2 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A4 = CLBLM_R_X15Y112_SLICE_X20Y112_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A5 = 1'b1;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_A6 = CLBLM_L_X16Y111_SLICE_X22Y111_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B1 = CLBLM_L_X16Y111_SLICE_X22Y111_DO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B3 = CLBLM_L_X16Y110_SLICE_X22Y110_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B4 = 1'b1;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B5 = CLBLM_R_X15Y112_SLICE_X20Y112_BO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_B6 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C1 = CLBLM_L_X16Y109_SLICE_X23Y109_AO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C2 = CLBLM_L_X16Y111_SLICE_X23Y111_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C3 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_C6 = CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D1 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D3 = CLBLM_L_X16Y111_SLICE_X23Y111_DO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D4 = CLBLM_L_X16Y109_SLICE_X22Y109_AO5;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_D6 = CLBLM_R_X15Y111_SLICE_X20Y111_AO6;
  assign CLBLM_L_X16Y111_SLICE_X22Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_R_X15Y116_SLICE_X20Y116_AQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLM_L_X16Y116_SLICE_X23Y116_BQ;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_D = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_D = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X15Y127_SLICE_X21Y127_B6 = CLBLM_R_X15Y127_SLICE_X21Y127_AO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A1 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A2 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A4 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_A6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B1 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B2 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B3 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B4 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_B6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C1 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C2 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C3 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C4 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_C6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D1 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D2 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D3 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D4 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X23Y113_D6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A2 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_A6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B1 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_B6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C2 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C3 = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_C6 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D1 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D2 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D3 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D4 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D5 = 1'b1;
  assign CLBLM_L_X16Y113_SLICE_X22Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = LIOB33_X0Y197_IOB_X0Y198_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y122_SLICE_X21Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A1 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A3 = CLBLM_L_X16Y114_SLICE_X22Y114_CO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A4 = CLBLM_L_X16Y115_SLICE_X23Y115_BQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_A6 = CLBLM_R_X15Y114_SLICE_X21Y114_BO5;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B1 = CLBLM_L_X16Y114_SLICE_X23Y114_DO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B3 = CLBLM_L_X16Y113_SLICE_X22Y113_AO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B4 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_B6 = CLBLM_L_X16Y114_SLICE_X22Y114_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B6 = 1'b1;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C1 = CLBLM_L_X16Y115_SLICE_X23Y115_BQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C3 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_C6 = CLBLM_L_X16Y113_SLICE_X22Y113_CO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A5 = CLBLM_R_X15Y122_SLICE_X20Y122_CO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_A6 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D1 = CLBLM_L_X16Y114_SLICE_X23Y114_BQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D3 = CLBLM_L_X16Y114_SLICE_X22Y114_BO5;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_D6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y114_SLICE_X23Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A1 = CLBLM_L_X16Y114_SLICE_X22Y114_DO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A4 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A5 = CLBLM_L_X16Y113_SLICE_X22Y113_BO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_A6 = CLBLM_R_X15Y114_SLICE_X21Y114_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B4 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B6 = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C1 = CLBLM_L_X16Y114_SLICE_X23Y114_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C5 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_C6 = CLBLM_L_X16Y113_SLICE_X22Y113_CO6;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D1 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D2 = CLBLM_L_X16Y114_SLICE_X22Y114_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D3 = CLBLM_L_X16Y113_SLICE_X22Y113_AO5;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_D6 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y114_SLICE_X22Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_L_X16Y117_SLICE_X22Y117_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D5 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D6 = CLBLM_R_X13Y124_SLICE_X18Y124_BQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_R_X15Y116_SLICE_X21Y116_BQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A4 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A6 = CLBLM_R_X13Y125_SLICE_X18Y125_CO6;
  assign CLBLM_L_X12Y123_SLICE_X17Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X15Y122_SLICE_X20Y122_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B6 = CLBLM_R_X15Y123_SLICE_X20Y123_BO6;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_D = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_D = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C2 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C4 = CLBLM_L_X16Y125_SLICE_X22Y125_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A1 = CLBLM_L_X16Y115_SLICE_X23Y115_DO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A2 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A4 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A5 = CLBLM_L_X16Y115_SLICE_X23Y115_CO5;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_A6 = CLBLM_L_X16Y115_SLICE_X22Y115_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B3 = CLBLM_L_X16Y115_SLICE_X23Y115_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B4 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B5 = CLBLM_L_X16Y114_SLICE_X23Y114_CO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_B6 = CLBLM_L_X16Y115_SLICE_X23Y115_CO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C3 = 1'b1;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C4 = CLBLM_R_X15Y115_SLICE_X21Y115_BO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C5 = 1'b1;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D2 = CLBLM_L_X16Y115_SLICE_X23Y115_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D3 = CLBLM_L_X16Y115_SLICE_X22Y115_DO6;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D4 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_D6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y115_SLICE_X23Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A1 = CLBLM_R_X15Y115_SLICE_X21Y115_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A3 = CLBLM_R_X15Y115_SLICE_X21Y115_BO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A5 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_A6 = CLBLM_L_X16Y115_SLICE_X22Y115_CO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B1 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B2 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B3 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B4 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_B6 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A6 = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C2 = CLBLM_L_X16Y115_SLICE_X22Y115_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C3 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C4 = CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C5 = CLBLM_L_X16Y116_SLICE_X23Y116_DO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_C6 = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D6 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D2 = 1'b1;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D4 = 1'b1;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D5 = 1'b1;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_D6 = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_L_X16Y115_SLICE_X22Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C1 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C2 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C5 = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_A6 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = CLBLM_R_X13Y122_SLICE_X18Y122_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A1 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A3 = CLBLM_L_X16Y114_SLICE_X23Y114_BQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A4 = CLBLM_L_X16Y114_SLICE_X22Y114_BO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_A6 = CLBLM_L_X16Y116_SLICE_X23Y116_CO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B1 = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B3 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B4 = CLBLM_L_X16Y116_SLICE_X22Y116_DO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_B6 = CLBLM_L_X16Y116_SLICE_X23Y116_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C2 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C4 = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C5 = CLBLM_L_X16Y116_SLICE_X23Y116_AQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_C6 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D2 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D4 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D5 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_D6 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X23Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A4 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A5 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B1 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B2 = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B4 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B5 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_B6 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C1 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C3 = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C5 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_C6 = 1'b1;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D2 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D3 = CLBLM_L_X16Y116_SLICE_X23Y116_DO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D4 = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D5 = CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  assign CLBLM_L_X16Y116_SLICE_X22Y116_D6 = CLBLM_L_X16Y116_SLICE_X23Y116_BQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A2 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A3 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A5 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_A6 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B2 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B3 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B4 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_B6 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C1 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C2 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C3 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C4 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C5 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_C6 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D1 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D2 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D3 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D4 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D5 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X19Y100_D6 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A2 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A3 = CLBLM_R_X13Y100_SLICE_X18Y100_BO5;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A4 = CLBLM_R_X13Y100_SLICE_X18Y100_DO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A5 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_A6 = CLBLM_R_X13Y104_SLICE_X18Y104_CO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B3 = CLBLM_L_X12Y101_SLICE_X17Y101_CO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B4 = CLBLM_R_X13Y100_SLICE_X18Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B5 = CLBLM_R_X15Y100_SLICE_X20Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_B6 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C1 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C2 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C3 = CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C4 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_C6 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLM_R_X15Y119_SLICE_X21Y119_BQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D1 = 1'b1;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D2 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D3 = CLBLM_R_X13Y100_SLICE_X19Y100_BO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D4 = CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X13Y100_SLICE_X18Y100_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_R_X15Y119_SLICE_X21Y119_AQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign RIOB33_X105Y101_IOB_X1Y102_O = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign RIOB33_X105Y101_IOB_X1Y101_O = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A1 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A2 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A3 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A4 = CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A5 = CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_A6 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B4 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_B6 = CLBLM_L_X16Y117_SLICE_X23Y117_AO5;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C1 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C2 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C3 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C4 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C5 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_C6 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D1 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D2 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D3 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D4 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D5 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X23Y117_D6 = 1'b1;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A2 = CLBLM_R_X15Y116_SLICE_X21Y116_BQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A4 = CLBLM_L_X16Y116_SLICE_X22Y116_BO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A5 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_A6 = CLBLM_L_X16Y117_SLICE_X22Y117_CO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B1 = CLBLM_L_X16Y117_SLICE_X22Y117_DO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B2 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B3 = CLBLM_L_X16Y117_SLICE_X22Y117_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_B6 = CLBLM_L_X16Y116_SLICE_X22Y116_AO5;
  assign LIOI3_X0Y147_ILOGIC_X0Y148_D = LIOB33_X0Y147_IOB_X0Y148_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_D = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C1 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C3 = CLBLM_L_X16Y117_SLICE_X22Y117_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C5 = CLBLM_L_X16Y116_SLICE_X22Y116_CO5;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_C6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D2 = CLBLM_L_X16Y116_SLICE_X22Y116_CO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D3 = CLBLM_L_X16Y117_SLICE_X22Y117_BQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D5 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_D6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y117_SLICE_X22Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A2 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A3 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A4 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A5 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_A6 = 1'b1;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B1 = CLBLM_R_X15Y101_SLICE_X21Y101_AO5;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B2 = CLBLM_R_X11Y102_SLICE_X15Y102_BO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B3 = CLBLM_R_X15Y100_SLICE_X20Y100_BO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B4 = CLBLM_R_X15Y101_SLICE_X20Y101_BO5;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B5 = CLBLM_R_X13Y101_SLICE_X19Y101_AO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_B6 = CLBLM_R_X13Y103_SLICE_X19Y103_CO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C1 = CLBLM_R_X13Y102_SLICE_X19Y102_AO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C2 = CLBLM_R_X13Y100_SLICE_X19Y100_BO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C3 = CLBLM_R_X13Y103_SLICE_X19Y103_AO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C4 = CLBLM_R_X15Y101_SLICE_X21Y101_BO5;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C5 = CLBLM_R_X15Y101_SLICE_X20Y101_AO5;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_C6 = CLBLM_R_X11Y101_SLICE_X15Y101_BO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D1 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D2 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D3 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D4 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D5 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_R_X13Y101_SLICE_X19Y101_D6 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A1 = CLBLM_R_X13Y103_SLICE_X18Y103_DO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A2 = CLBLM_R_X13Y101_SLICE_X18Y101_DO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A3 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A5 = 1'b1;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_A6 = CLBLM_R_X13Y101_SLICE_X18Y101_CO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B2 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B3 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B4 = CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_B6 = 1'b1;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C1 = CLBLM_R_X13Y102_SLICE_X19Y102_AO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C2 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C5 = CLBLM_R_X13Y101_SLICE_X18Y101_BO5;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_C6 = 1'b1;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D1 = 1'b1;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D2 = CLBLM_R_X13Y101_SLICE_X19Y101_AO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D5 = 1'b1;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_D6 = CLBLM_L_X12Y102_SLICE_X17Y102_BO6;
  assign CLBLM_R_X13Y101_SLICE_X18Y101_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y103_IOB_X1Y104_O = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign RIOB33_X105Y103_IOB_X1Y103_O = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A4 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A1 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A2 = CLBLM_R_X15Y117_SLICE_X21Y117_BQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A3 = CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A4 = CLBLM_L_X16Y118_SLICE_X23Y118_BO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B3 = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B4 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_B6 = CLBLM_L_X16Y118_SLICE_X23Y118_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C1 = CLBLM_R_X15Y115_SLICE_X21Y115_DO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C2 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C3 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C4 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C5 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_C6 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D1 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D2 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D3 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D4 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D5 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A6 = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_L_X16Y118_SLICE_X23Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A1 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A2 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A3 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A4 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A5 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_A6 = CLBLM_R_X15Y118_SLICE_X20Y118_DO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B2 = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B1 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B2 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B3 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B4 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B5 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B3 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B4 = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C1 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C2 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C3 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C4 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C5 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_C6 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D1 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D2 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D3 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D4 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D5 = 1'b1;
  assign CLBLM_L_X16Y118_SLICE_X22Y118_D6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A1 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A2 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A3 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A4 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A5 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_A6 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B2 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B3 = CLBLM_L_X12Y102_SLICE_X17Y102_DO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B4 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B5 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_B6 = CLBLM_R_X13Y102_SLICE_X19Y102_AO5;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C2 = CLBLM_L_X12Y102_SLICE_X17Y102_DO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C4 = CLBLM_R_X13Y102_SLICE_X19Y102_AO5;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C5 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D1 = CLBLM_R_X15Y102_SLICE_X21Y102_AO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D2 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D4 = CLBLM_R_X13Y102_SLICE_X19Y102_CO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X13Y102_SLICE_X19Y102_D6 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A2 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A3 = CLBLM_R_X13Y103_SLICE_X19Y103_DO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A4 = CLBLM_R_X13Y102_SLICE_X18Y102_BO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A5 = CLBLM_R_X13Y102_SLICE_X18Y102_CO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_A6 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B1 = CLBLM_R_X13Y103_SLICE_X19Y103_CO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B2 = CLBLM_R_X13Y103_SLICE_X18Y103_BO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B3 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B5 = CLBLM_R_X13Y101_SLICE_X18Y101_BO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_B6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign RIOB33_X105Y105_IOB_X1Y106_O = CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  assign RIOB33_X105Y105_IOB_X1Y105_O = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C1 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C2 = CLBLM_L_X12Y103_SLICE_X17Y103_CO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C5 = CLBLM_R_X13Y103_SLICE_X19Y103_CO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_C6 = CLBLM_R_X13Y103_SLICE_X19Y103_AO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D1 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D2 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D3 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D4 = CLBLM_L_X12Y102_SLICE_X17Y102_DO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D5 = 1'b1;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_D6 = CLBLM_R_X13Y103_SLICE_X19Y103_AO6;
  assign CLBLM_R_X13Y102_SLICE_X18Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A6 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X15Y123_SLICE_X21Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A1 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A4 = CLBLM_L_X16Y119_SLICE_X23Y119_BO6;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A5 = CLBLM_L_X16Y119_SLICE_X22Y119_BO5;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_A6 = CLBLM_R_X15Y119_SLICE_X20Y119_AQ;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B3 = CLBLM_L_X16Y119_SLICE_X23Y119_AQ;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B5 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_B6 = CLBLM_R_X15Y119_SLICE_X20Y119_BO6;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C1 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C2 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C3 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C4 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C5 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_C6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A5 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D1 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D2 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D3 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D4 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D5 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_D6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A5 = CLBLM_R_X15Y123_SLICE_X20Y123_CO5;
  assign CLBLM_L_X16Y119_SLICE_X23Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A1 = CLBLM_L_X16Y119_SLICE_X22Y119_DO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A2 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A3 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A4 = CLBLM_L_X16Y119_SLICE_X22Y119_BO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A5 = CLBLM_L_X16Y119_SLICE_X23Y119_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B2 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B1 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B2 = CLBLM_R_X15Y117_SLICE_X21Y117_CO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B3 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B4 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B5 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_B6 = 1'b1;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C1 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C2 = CLBLM_R_X15Y118_SLICE_X20Y118_DO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C3 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C4 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C5 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B5 = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B6 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D1 = CLBLM_L_X16Y119_SLICE_X22Y119_CO5;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D2 = CLBLM_L_X16Y119_SLICE_X22Y119_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D5 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X16Y119_SLICE_X22Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C4 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A1 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A3 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A4 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A5 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B1 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B3 = CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B4 = CLBLM_L_X12Y103_SLICE_X17Y103_CO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B5 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_B6 = CLBLM_R_X13Y103_SLICE_X19Y103_CO6;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C3 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C4 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_C6 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D2 = CLBLM_R_X13Y102_SLICE_X18Y102_DO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D3 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D6 = 1'b1;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D5 = CLBLM_R_X15Y108_SLICE_X20Y108_BO6;
  assign CLBLM_R_X13Y103_SLICE_X19Y103_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign RIOB33_X105Y107_IOB_X1Y107_O = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign RIOB33_X105Y107_IOB_X1Y108_O = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A1 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A2 = CLBLM_R_X13Y103_SLICE_X19Y103_BO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A3 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A4 = CLBLM_R_X13Y103_SLICE_X18Y103_BO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_A6 = CLBLM_R_X13Y102_SLICE_X18Y102_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B4 = CLBLM_L_X12Y103_SLICE_X17Y103_BO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B5 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_B6 = 1'b1;
  assign CLBLM_R_X15Y123_SLICE_X20Y123_D6 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C1 = CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C4 = CLBLM_L_X12Y102_SLICE_X17Y102_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C5 = CLBLM_R_X15Y108_SLICE_X20Y108_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_C6 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D3 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D4 = CLBLM_L_X12Y102_SLICE_X17Y102_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D5 = CLBLM_R_X15Y108_SLICE_X20Y108_CO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_D6 = CLBLM_L_X12Y103_SLICE_X17Y103_DO6;
  assign CLBLM_R_X13Y103_SLICE_X18Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C5 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A1 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A2 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A3 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A4 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A5 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_A6 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B1 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B2 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B3 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B4 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B5 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_B6 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C1 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C2 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C3 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C4 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C5 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_C6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D1 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D2 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D3 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D4 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D5 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X13Y100_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A4 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A5 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D6 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B1 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B2 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B3 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B4 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B5 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_B6 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C1 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C4 = CLBLM_L_X10Y100_SLICE_X12Y100_AO5;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C5 = CLBLM_L_X10Y101_SLICE_X13Y101_AO5;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_C6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D1 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D2 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D3 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D4 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D5 = 1'b1;
  assign CLBLM_L_X10Y100_SLICE_X12Y100_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A1 = CLBLM_R_X13Y102_SLICE_X19Y102_DO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A2 = CLBLM_R_X15Y102_SLICE_X20Y102_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C2 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A5 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_A6 = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C3 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign RIOB33_X105Y109_IOB_X1Y109_O = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B1 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B2 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B3 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B4 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B5 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_B6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C1 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C2 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C6 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C3 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C4 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C5 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_C6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D1 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D2 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D3 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D4 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D5 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_D6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X19Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A2 = CLBLM_R_X13Y100_SLICE_X18Y100_BO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A3 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A4 = CLBLM_R_X13Y104_SLICE_X18Y104_BO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_A6 = CLBLM_R_X13Y103_SLICE_X18Y103_BO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B1 = CLBLM_R_X13Y104_SLICE_X18Y104_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C4 = CLBLM_R_X13Y103_SLICE_X18Y103_BO5;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C5 = CLBLM_R_X13Y104_SLICE_X18Y104_DO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_C6 = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D1 = CLBLM_L_X12Y101_SLICE_X17Y101_AO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D2 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D4 = CLBLM_R_X13Y100_SLICE_X19Y100_BO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D5 = 1'b1;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_D6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X13Y104_SLICE_X18Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_A6 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B3 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X23Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A2 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A4 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A5 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A6 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A1 = CLBLM_R_X15Y122_SLICE_X20Y122_AQ;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A2 = CLBLM_L_X16Y123_SLICE_X22Y123_AO6;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A3 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A5 = CLBLM_R_X15Y121_SLICE_X21Y121_BO6;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_A6 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B1 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B2 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C1 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C2 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D1 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D3 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D4 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D5 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D6 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D1 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D2 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D3 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D4 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D5 = 1'b1;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A1 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A2 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A3 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X16Y121_SLICE_X22Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A4 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A5 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B2 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B3 = CLBLM_L_X10Y100_SLICE_X12Y100_AO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B5 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B6 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C1 = CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C2 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C3 = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C6 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D1 = CLBLM_R_X11Y100_SLICE_X14Y100_AO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D2 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D3 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D4 = CLBLM_L_X10Y101_SLICE_X12Y101_AO5;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D5 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D6 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  assign RIOB33_X105Y111_IOB_X1Y111_O = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = LIOB33_X0Y183_IOB_X0Y184_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = LIOB33_X0Y183_IOB_X0Y184_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = 1'b1;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A1 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A2 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A3 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A4 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A5 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A6 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B1 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B2 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B3 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B4 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B5 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B6 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C1 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C2 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C3 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C4 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C5 = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C6 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D6 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A1 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A2 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A4 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A5 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B1 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B3 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B4 = CLBLM_L_X10Y100_SLICE_X12Y100_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B6 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign LIOI3_SING_X0Y149_ILOGIC_X0Y149_D = LIOB33_SING_X0Y149_IOB_X0Y149_I;
  assign RIOB33_X105Y113_IOB_X1Y114_O = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C1 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C2 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C3 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C5 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C6 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D4 = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D6 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A1 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A2 = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A3 = CLBLM_R_X15Y108_SLICE_X20Y108_BO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A5 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A6 = CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D6 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A1 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A2 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A3 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A4 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A5 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A6 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B4 = CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B3 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B5 = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B6 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C2 = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C3 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C6 = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D2 = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D3 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D4 = CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C1 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C2 = CLBLM_R_X13Y103_SLICE_X19Y103_AO5;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A1 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A2 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A3 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A4 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A5 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_A6 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B1 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B2 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B3 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B4 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B5 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_B6 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C1 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C2 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C3 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C4 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C5 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_C6 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D1 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D2 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D3 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D4 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D5 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X23Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A1 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A2 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A5 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A6 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B2 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B2 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_B6 = CLBLM_R_X15Y124_SLICE_X21Y124_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C1 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C2 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C1 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C2 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C3 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C4 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C5 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_C6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D1 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D2 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D5 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D6 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign RIOB33_X105Y115_IOB_X1Y115_O = CLBLM_R_X15Y114_SLICE_X21Y114_AQ;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D1 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D2 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D3 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D4 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D5 = 1'b1;
  assign CLBLM_L_X16Y123_SLICE_X22Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A1 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A2 = CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A3 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A5 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B1 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B2 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B3 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B5 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B6 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C1 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C2 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C3 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C5 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C6 = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D2 = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D6 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A1 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A2 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A3 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A4 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A5 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B1 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B2 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B3 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B4 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B5 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B6 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C1 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C2 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C3 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C4 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C5 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C6 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D1 = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D2 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D3 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D6 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C4 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C5 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C6 = 1'b1;
  assign CLBLM_R_X15Y124_SLICE_X21Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A3 = CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A4 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A5 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A6 = CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLM_L_X16Y116_SLICE_X23Y116_AQ;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A5 = CLBLM_R_X15Y124_SLICE_X20Y124_CO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B1 = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B2 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B3 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B5 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_A6 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign RIOB33_X105Y117_IOB_X1Y117_O = CLBLM_L_X16Y114_SLICE_X23Y114_BQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C1 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C5 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C6 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D1 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D3 = CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D5 = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A3 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A4 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A5 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A6 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B2 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B5 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B6 = 1'b1;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y124_SLICE_X20Y124_B6 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C1 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C3 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C4 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D2 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D3 = CLBLM_L_X10Y102_SLICE_X12Y102_BQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D4 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D5 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D6 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A1 = CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A2 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A4 = CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A5 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B1 = CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B2 = CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B3 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B5 = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B6 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C1 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C2 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C3 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C4 = CLBLM_R_X13Y108_SLICE_X19Y108_AO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C5 = CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C6 = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D1 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D3 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D6 = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A2 = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A3 = CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A5 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B1 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B2 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B3 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B4 = CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B5 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B6 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A6 = CLBLM_R_X13Y126_SLICE_X18Y126_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C1 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C2 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C3 = CLBLM_R_X13Y103_SLICE_X18Y103_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C4 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C5 = CLBLM_R_X13Y104_SLICE_X18Y104_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C6 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D4 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C1 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C2 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B1 = CLBLM_R_X15Y127_SLICE_X21Y127_AO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B2 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B3 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B4 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B5 = CLBLM_L_X16Y125_SLICE_X23Y125_AO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_R_X15Y116_SLICE_X20Y116_AQ;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLM_L_X16Y116_SLICE_X23Y116_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C5 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C2 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C3 = CLBLM_L_X16Y125_SLICE_X23Y125_AO5;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C4 = CLBLM_R_X15Y127_SLICE_X21Y127_AO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_C6 = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C6 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_D = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D1 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D3 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D5 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X16Y125_SLICE_X23Y125_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_D = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A1 = CLBLM_L_X16Y126_SLICE_X22Y126_AQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A2 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A4 = CLBLM_L_X16Y125_SLICE_X22Y125_BO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A5 = CLBLM_L_X16Y125_SLICE_X22Y125_CO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_A6 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_B6 = 1'b1;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C2 = CLBLM_L_X16Y125_SLICE_X22Y125_AQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C3 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C5 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D2 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D3 = CLBLM_L_X16Y125_SLICE_X23Y125_DO6;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_L_X16Y125_SLICE_X22Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D6 = CLBLM_L_X16Y125_SLICE_X23Y125_CO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A3 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A6 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B2 = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B3 = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A2 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A3 = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A4 = CLBLM_R_X15Y108_SLICE_X20Y108_AO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A5 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A6 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B2 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B3 = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B5 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B6 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C1 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C2 = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C6 = CLBLM_R_X15Y108_SLICE_X20Y108_AO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D3 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D6 = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLM_R_X15Y115_SLICE_X20Y115_AQ;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLM_R_X15Y116_SLICE_X20Y116_BQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A2 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_A6 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B2 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_B6 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C1 = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C2 = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C4 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_C6 = CLBLM_L_X16Y125_SLICE_X23Y125_AO5;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D1 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D2 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D3 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D4 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X16Y126_SLICE_X23Y126_D6 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A6 = CLBLM_L_X16Y126_SLICE_X22Y126_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B6 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C2 = CLBLM_L_X16Y126_SLICE_X22Y126_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = 1'b1;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C3 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C4 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C6 = 1'b1;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D6 = 1'b1;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A1 = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A2 = CLBLM_R_X15Y110_SLICE_X20Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A3 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A6 = CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B1 = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B3 = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B4 = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B6 = CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C1 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C2 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C4 = CLBLM_L_X16Y109_SLICE_X23Y109_AO5;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C5 = CLBLM_R_X13Y112_SLICE_X18Y112_BO5;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C6 = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D1 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D6 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLM_L_X16Y115_SLICE_X22Y115_AQ;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLM_R_X15Y115_SLICE_X21Y115_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = CLBLM_L_X8Y103_SLICE_X11Y103_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A3 = CLBLM_L_X16Y109_SLICE_X22Y109_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B1 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B5 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_B6 = CLBLM_R_X13Y111_SLICE_X19Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C2 = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C3 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C4 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_C6 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D1 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D2 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D3 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D4 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D5 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X19Y111_D6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A1 = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A4 = CLBLM_R_X13Y111_SLICE_X18Y111_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A5 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_A6 = CLBLM_R_X13Y114_SLICE_X18Y114_BO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B3 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B5 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_B6 = 1'b1;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C1 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C2 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C3 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C5 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_C6 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_L_X16Y115_SLICE_X23Y115_AQ;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLM_L_X16Y115_SLICE_X23Y115_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D2 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D3 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_D6 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_R_X13Y111_SLICE_X18Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C1 = CLBLM_R_X15Y100_SLICE_X21Y100_AO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C2 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A4 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y125_SLICE_X21Y125_A6 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A1 = CLBLM_L_X16Y109_SLICE_X22Y109_DO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B1 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B4 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B5 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B6 = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C1 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C2 = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C3 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C4 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C5 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D6 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_L_X16Y114_SLICE_X23Y114_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A1 = CLBLM_R_X15Y107_SLICE_X21Y107_CQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B1 = CLBLM_L_X12Y115_SLICE_X16Y115_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B3 = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B4 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C1 = CLBLM_L_X16Y109_SLICE_X23Y109_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C3 = CLBLM_R_X15Y110_SLICE_X21Y110_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C4 = CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C5 = CLBLM_L_X16Y109_SLICE_X22Y109_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C6 = CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D1 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D2 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D3 = CLBLM_R_X15Y112_SLICE_X20Y112_AO5;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D4 = CLBLM_L_X12Y115_SLICE_X16Y115_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A2 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A3 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A4 = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A5 = CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B1 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B6 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_R_X15Y114_SLICE_X20Y114_AQ;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_R_X15Y116_SLICE_X21Y116_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C1 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C2 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C3 = CLBLM_R_X13Y114_SLICE_X18Y114_AO5;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C4 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C5 = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C6 = CLBLM_R_X15Y110_SLICE_X20Y110_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D1 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D2 = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D4 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D5 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A1 = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A2 = CLBLM_R_X15Y110_SLICE_X20Y110_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A4 = CLBLM_R_X13Y114_SLICE_X18Y114_AO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A5 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A6 = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B1 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B3 = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B6 = CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C1 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C2 = CLBLM_R_X15Y112_SLICE_X20Y112_AO5;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C3 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C5 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C6 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A6 = CLBLM_R_X13Y130_SLICE_X18Y130_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D1 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D2 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D3 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D4 = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D5 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B6 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A6 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_L_X16Y117_SLICE_X22Y117_AQ;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_R_X15Y116_SLICE_X21Y116_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A1 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A3 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A4 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A5 = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_A6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C1 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_C6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D1 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C5 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D3 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D4 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C6 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X13Y114_SLICE_X19Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A1 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A2 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A4 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A5 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_A6 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B1 = CLBLM_R_X13Y114_SLICE_X18Y114_DO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B2 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B4 = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B5 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_B6 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C1 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C2 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C3 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C4 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C5 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_C6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D1 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D2 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D3 = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D4 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D5 = 1'b1;
  assign CLBLM_R_X13Y114_SLICE_X18Y114_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D3 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_L_X16Y117_SLICE_X22Y117_BQ;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_R_X15Y117_SLICE_X21Y117_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_A6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_B6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_C6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D1 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D2 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D3 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D4 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D5 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X19Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A1 = CLBLM_L_X16Y115_SLICE_X22Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A2 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A3 = CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A4 = CLBLM_R_X13Y115_SLICE_X18Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_A6 = 1'b1;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B1 = CLBLM_R_X13Y115_SLICE_X18Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B4 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_B6 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C2 = CLBLM_L_X12Y116_SLICE_X16Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C3 = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C4 = CLBLM_L_X12Y116_SLICE_X16Y116_A5Q;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C5 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_C6 = CLBLM_L_X12Y116_SLICE_X17Y116_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D1 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D2 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D4 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D5 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_D6 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_R_X13Y115_SLICE_X18Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B3 = CLBLM_R_X15Y103_SLICE_X20Y103_AO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B4 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C1 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C2 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_R_X15Y117_SLICE_X21Y117_AQ;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_R_X15Y117_SLICE_X20Y117_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D5 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D6 = CLBLM_R_X15Y106_SLICE_X20Y106_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A1 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A3 = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A4 = CLBLM_L_X16Y117_SLICE_X23Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A5 = CLBLM_R_X13Y115_SLICE_X18Y115_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A6 = CLBLM_R_X13Y115_SLICE_X18Y115_AO5;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B5 = CLBLM_L_X10Y103_SLICE_X12Y103_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B6 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C4 = CLBLM_L_X8Y102_SLICE_X11Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C5 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C6 = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLM_R_X15Y119_SLICE_X20Y119_AQ;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLM_R_X15Y118_SLICE_X20Y118_AQ;
  assign CLBLM_R_X15Y126_SLICE_X21Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = CLBLM_R_X11Y114_SLICE_X15Y114_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A5 = CLBLM_L_X16Y126_SLICE_X22Y126_BO5;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_A6 = CLBLM_R_X15Y126_SLICE_X20Y126_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_L_X10Y114_SLICE_X12Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C2 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A6 = 1'b1;
  assign CLBLM_R_X15Y126_SLICE_X20Y126_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D6 = 1'b1;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_L_X16Y119_SLICE_X22Y119_AQ;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_L_X16Y119_SLICE_X23Y119_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C1 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C5 = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_AX = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_BX = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D6 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y122_SLICE_X16Y122_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A1 = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A2 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A6 = CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D3 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D5 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D6 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLM_R_X15Y119_SLICE_X21Y119_BQ;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_R_X15Y119_SLICE_X21Y119_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_D = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_AX = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A1 = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A2 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A3 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A5 = CLBLM_R_X15Y122_SLICE_X21Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A6 = CLBLM_R_X13Y121_SLICE_X19Y121_BO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B2 = CLBLM_R_X15Y121_SLICE_X20Y121_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B3 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B5 = CLBLM_R_X15Y122_SLICE_X21Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B6 = CLBLM_R_X15Y122_SLICE_X20Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C6 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D1 = CLBLM_R_X15Y122_SLICE_X21Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D2 = CLBLM_R_X15Y121_SLICE_X20Y121_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D4 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D5 = CLBLM_R_X15Y122_SLICE_X20Y122_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A3 = CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A6 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B3 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B4 = CLBLM_L_X16Y121_SLICE_X22Y121_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B5 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B6 = CLBLM_R_X15Y120_SLICE_X20Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C2 = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C3 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C6 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLM_R_X15Y132_SLICE_X21Y132_AQ;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLM_R_X15Y118_SLICE_X21Y118_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D1 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D2 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D4 = CLBLM_R_X15Y120_SLICE_X20Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D6 = CLBLM_L_X16Y121_SLICE_X22Y121_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A1 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A3 = 1'b1;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A5 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_A6 = CLBLM_R_X13Y121_SLICE_X19Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B3 = CLBLM_R_X13Y120_SLICE_X19Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B4 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C2 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C3 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C5 = CLBLM_R_X13Y121_SLICE_X19Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_C6 = CLBLM_R_X13Y121_SLICE_X19Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D5 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y121_SLICE_X19Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_R_X15Y132_SLICE_X21Y132_CQ;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLM_R_X15Y132_SLICE_X21Y132_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A1 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A3 = CLBLM_R_X13Y125_SLICE_X18Y125_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A4 = CLBLM_R_X15Y121_SLICE_X20Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_A6 = CLBLM_R_X13Y121_SLICE_X18Y121_CO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B2 = CLBLM_R_X15Y121_SLICE_X21Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B3 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B4 = CLBLM_R_X15Y121_SLICE_X20Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_B6 = CLBLM_R_X15Y120_SLICE_X21Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C2 = CLBLM_R_X13Y121_SLICE_X18Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C3 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C4 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_C6 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D1 = CLBLM_L_X12Y120_SLICE_X16Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D2 = CLBLM_R_X15Y121_SLICE_X21Y121_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D4 = CLBLM_R_X15Y121_SLICE_X20Y121_BQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_D6 = CLBLM_R_X15Y120_SLICE_X21Y120_AQ;
  assign CLBLM_R_X13Y121_SLICE_X18Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A1 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A2 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A5 = CLBLM_R_X13Y124_SLICE_X19Y124_BO5;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_A6 = CLBLM_R_X13Y122_SLICE_X19Y122_CO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B1 = CLBLM_R_X15Y122_SLICE_X20Y122_BQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B3 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B4 = CLBLM_R_X15Y123_SLICE_X21Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_B6 = CLBLM_R_X15Y123_SLICE_X20Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C1 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C2 = CLBLM_L_X16Y125_SLICE_X23Y125_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C5 = CLBLM_R_X13Y122_SLICE_X19Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D1 = CLBLM_L_X12Y122_SLICE_X16Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D2 = CLBLM_R_X15Y123_SLICE_X20Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D5 = CLBLM_R_X15Y122_SLICE_X20Y122_BQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A3 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A4 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A5 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A6 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_D6 = CLBLM_R_X15Y123_SLICE_X21Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A1 = CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B3 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B5 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B6 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A2 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A3 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A4 = CLBLM_R_X13Y122_SLICE_X18Y122_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C2 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B3 = CLBLM_R_X13Y122_SLICE_X18Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B4 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D2 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C3 = CLBLM_L_X12Y123_SLICE_X17Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C4 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A2 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D3 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D4 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D5 = CLBLM_L_X12Y122_SLICE_X17Y122_AQ;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B2 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B6 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C2 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D2 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A1 = CLBLM_R_X13Y123_SLICE_X19Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A3 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A4 = CLBLM_R_X13Y123_SLICE_X19Y123_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A5 = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C5 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D1 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D3 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D4 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D5 = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A2 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A3 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A5 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_D6 = CLBLM_L_X12Y123_SLICE_X17Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A1 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B3 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A2 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_A4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C1 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C2 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C5 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C6 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B1 = CLBLM_R_X13Y123_SLICE_X18Y123_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B3 = CLBLM_R_X13Y123_SLICE_X18Y123_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B4 = CLBLM_R_X13Y123_SLICE_X19Y123_CO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B5 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D1 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D3 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D5 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D6 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C4 = CLBLM_R_X15Y127_SLICE_X21Y127_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D3 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D4 = CLBLM_R_X13Y123_SLICE_X18Y123_BQ;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_D5 = CLBLM_L_X16Y125_SLICE_X22Y125_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B1 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X18Y123_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y127_SLICE_X20Y127_D6 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C1 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C2 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C3 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C5 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C6 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D1 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D3 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D4 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D5 = CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C2 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C5 = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C6 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = CLBLM_L_X16Y111_SLICE_X23Y111_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A4 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A5 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_A6 = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A1 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A2 = CLBLM_R_X15Y124_SLICE_X20Y124_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A4 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A5 = CLBLM_L_X16Y125_SLICE_X22Y125_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_A6 = CLBLM_R_X13Y124_SLICE_X19Y124_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C1 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C3 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_C6 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D1 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D3 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X13Y124_SLICE_X19Y124_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A5 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_B6 = CLBLM_L_X16Y123_SLICE_X22Y123_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B3 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B5 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A2 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_A3 = CLBLM_L_X16Y123_SLICE_X22Y123_AO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C1 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C2 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C3 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C4 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C5 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C6 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B1 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B3 = CLBLM_R_X13Y124_SLICE_X19Y124_DO6;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B4 = CLBLM_R_X13Y127_SLICE_X19Y127_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D1 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D2 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D3 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D5 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D6 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_C6 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A1 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A6 = 1'b1;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D2 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X13Y124_SLICE_X18Y124_D4 = CLBLM_L_X16Y125_SLICE_X22Y125_AQ;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B3 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_C6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B4 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B5 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B6 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C1 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C2 = CLBLM_L_X8Y102_SLICE_X10Y102_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C3 = CLBLM_L_X8Y103_SLICE_X10Y103_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C4 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C5 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C6 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_L_X12Y123_SLICE_X16Y123_D6 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = CLBLM_R_X15Y125_SLICE_X20Y125_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = CLBLM_R_X13Y122_SLICE_X19Y122_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A2 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A3 = CLBLM_R_X13Y124_SLICE_X19Y124_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A4 = CLBLM_R_X15Y125_SLICE_X20Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_A5 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B2 = CLBLM_R_X15Y125_SLICE_X21Y125_BQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B4 = CLBLM_R_X13Y130_SLICE_X18Y130_BQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B5 = CLBLM_R_X15Y124_SLICE_X20Y124_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_B6 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C1 = CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C2 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C4 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C5 = CLBLM_R_X13Y125_SLICE_X19Y125_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D1 = CLBLM_R_X15Y124_SLICE_X20Y124_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D2 = CLBLM_R_X15Y125_SLICE_X21Y125_BQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X19Y125_D6 = CLBLM_R_X13Y130_SLICE_X18Y130_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A1 = CLBLM_R_X13Y125_SLICE_X18Y125_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A2 = CLBLM_R_X13Y124_SLICE_X18Y124_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A3 = CLBLM_R_X15Y125_SLICE_X21Y125_CO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_A4 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C3 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_C6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = 1'b1;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D3 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_D5 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X13Y125_SLICE_X18Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = CLBLM_R_X15Y125_SLICE_X20Y125_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_R_X13Y122_SLICE_X19Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = CLBLM_R_X15Y125_SLICE_X20Y125_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLM_R_X13Y124_SLICE_X18Y124_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = CLBLM_R_X13Y124_SLICE_X18Y124_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = CLBLM_R_X13Y122_SLICE_X18Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A1 = CLBLM_R_X13Y126_SLICE_X19Y126_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A2 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A5 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_A6 = CLBLM_R_X15Y122_SLICE_X20Y122_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B1 = CLBLM_L_X16Y125_SLICE_X22Y125_BO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B3 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B4 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B5 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_B6 = CLBLM_R_X13Y126_SLICE_X19Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C1 = CLBLM_R_X13Y126_SLICE_X19Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C2 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C4 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_C6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D3 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D4 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y126_SLICE_X19Y126_D6 = CLBLM_R_X13Y126_SLICE_X19Y126_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A1 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A3 = CLBLM_R_X15Y125_SLICE_X21Y125_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_A4 = CLBLM_R_X13Y125_SLICE_X18Y125_BO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B1 = CLBLM_R_X13Y126_SLICE_X18Y126_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B2 = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B3 = CLBLM_L_X12Y124_SLICE_X17Y124_AQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B4 = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C3 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = 1'b1;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D3 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D4 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_D5 = CLBLM_R_X15Y126_SLICE_X21Y126_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X13Y126_SLICE_X18Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = CLBLM_R_X13Y127_SLICE_X19Y127_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = CLBLM_R_X13Y127_SLICE_X19Y127_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_D = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = CLBLM_L_X12Y122_SLICE_X16Y122_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = CLBLM_R_X13Y125_SLICE_X19Y125_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = CLBLM_L_X12Y122_SLICE_X16Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = CLBLM_L_X12Y125_SLICE_X17Y125_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A1 = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A2 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A4 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A5 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A6 = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B2 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B3 = CLBLM_L_X12Y127_SLICE_X17Y127_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B4 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B5 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B6 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D1 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D2 = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D4 = CLBLM_R_X13Y127_SLICE_X19Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = LIOB33_X0Y147_IOB_X0Y148_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D6 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B1 = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B2 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B4 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B5 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = 1'b1;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y101_SLICE_X22Y101_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = CLBLM_L_X12Y124_SLICE_X17Y124_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = CLBLM_R_X11Y127_SLICE_X14Y127_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A2 = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A3 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A4 = CLBLM_R_X15Y120_SLICE_X21Y120_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A6 = CLBLM_R_X15Y128_SLICE_X20Y128_BO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B2 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B4 = CLBLM_L_X16Y126_SLICE_X23Y126_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C1 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C3 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C4 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C5 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C6 = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D1 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D2 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D4 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B2 = CLBLM_L_X12Y127_SLICE_X16Y127_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B3 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B5 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B6 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C3 = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C4 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C6 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A6 = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D6 = CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_A5Q;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_T1 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C2 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_T1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C5 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = CLBLM_R_X15Y125_SLICE_X20Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = CLBLM_R_X15Y130_SLICE_X20Y130_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D6 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A4 = CLBLM_L_X12Y124_SLICE_X16Y124_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A1 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_A6 = CLBLM_R_X15Y127_SLICE_X21Y127_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A2 = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A4 = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A5 = CLBLM_L_X12Y127_SLICE_X17Y127_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A6 = 1'b1;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_D = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_D = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B1 = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B2 = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B3 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B4 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B6 = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D2 = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D6 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B1 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B2 = CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B5 = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B6 = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C3 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C4 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_C5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D3 = CLBLM_R_X13Y124_SLICE_X19Y124_AQ;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D5 = CLBLM_R_X13Y125_SLICE_X18Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X12Y124_SLICE_X16Y124_D6 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = CLBLM_R_X13Y126_SLICE_X18Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = CLBLM_R_X11Y130_SLICE_X15Y130_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A1 = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A3 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A4 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A6 = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C2 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C3 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C4 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C5 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C6 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A2 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A4 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B1 = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B3 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B4 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C3 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C4 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C6 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D1 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D2 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D3 = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D4 = CLBLM_R_X13Y130_SLICE_X18Y130_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D5 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = CLBLM_R_X11Y131_SLICE_X14Y131_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_D1 = CLBLM_L_X10Y119_SLICE_X13Y119_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_D1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A2 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B1 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B2 = CLBLM_R_X15Y126_SLICE_X20Y126_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B5 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B6 = CLBLM_R_X15Y126_SLICE_X21Y126_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C2 = CLBLM_R_X15Y126_SLICE_X21Y126_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C3 = CLBLM_R_X15Y126_SLICE_X20Y126_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C4 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C5 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D2 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D3 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D4 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A1 = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A4 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B2 = CLBLM_R_X15Y130_SLICE_X20Y130_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C1 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C2 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C3 = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C4 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C5 = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D2 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D3 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D5 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_A5Q;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = 1'b1;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_D = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_D = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = CLBLM_R_X13Y126_SLICE_X18Y126_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = CLBLM_L_X16Y126_SLICE_X23Y126_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = CLBLM_L_X16Y126_SLICE_X23Y126_AO5;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = CLBLM_R_X11Y129_SLICE_X15Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A5 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B4 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C1 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C2 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C4 = CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C5 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C6 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B1 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B2 = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B3 = CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B5 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C3 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = 1'b1;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X16Y102_SLICE_X22Y102_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_C5 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_R_X13Y122_SLICE_X19Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = CLBLM_L_X12Y129_SLICE_X16Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_R_X15Y117_SLICE_X20Y117_AQ;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A6 = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_R_X15Y117_SLICE_X21Y117_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B5 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B6 = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_A6 = CLBLM_R_X13Y123_SLICE_X19Y123_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = CLBLM_R_X11Y125_SLICE_X15Y125_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = CLBLM_L_X10Y130_SLICE_X13Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_D = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_D = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D6 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_A6 = CLBLM_L_X12Y125_SLICE_X16Y125_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_L_X12Y115_SLICE_X17Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C2 = CLBLM_L_X12Y125_SLICE_X16Y125_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y120_SLICE_X20Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  assign CLBLM_L_X12Y125_SLICE_X16Y125_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = CLBLM_R_X11Y129_SLICE_X15Y129_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = CLBLM_L_X8Y130_SLICE_X11Y130_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X13Y122_SLICE_X18Y122_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = CLBLM_R_X15Y107_SLICE_X21Y107_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = CLBLM_R_X15Y127_SLICE_X21Y127_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = CLBLM_R_X13Y114_SLICE_X19Y114_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = CLBLM_R_X13Y111_SLICE_X18Y111_BO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_D = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_D = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = 1'b1;
  assign CLBLM_L_X16Y103_SLICE_X22Y103_B6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_B5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A6 = CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = CLBLM_L_X16Y114_SLICE_X22Y114_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = CLBLM_R_X15Y114_SLICE_X21Y114_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C2 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y116_SLICE_X0Y116_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C5 = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D6 = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_D = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_D = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B6 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A4 = CLBLM_L_X16Y126_SLICE_X22Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y115_SLICE_X0Y115_B5Q;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A6 = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C1 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C5 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C6 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLM_L_X16Y116_SLICE_X23Y116_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = CLBLM_L_X16Y114_SLICE_X23Y114_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_D = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_D = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A1 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A2 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A3 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A4 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A5 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_A6 = CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B1 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B2 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B3 = CLBLM_L_X12Y101_SLICE_X17Y101_CO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B4 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B5 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_B6 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C1 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C2 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C4 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C5 = CLBLM_L_X12Y101_SLICE_X17Y101_CO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_C6 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B3 = CLBLM_L_X16Y104_SLICE_X22Y104_DO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B4 = CLBLM_R_X15Y105_SLICE_X20Y105_DO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D1 = CLBLM_L_X12Y100_SLICE_X17Y100_AO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D2 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D3 = CLBLM_R_X15Y100_SLICE_X20Y100_BO5;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B5 = CLBLM_L_X16Y103_SLICE_X22Y103_AO6;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D5 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y100_SLICE_X21Y100_D6 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_B6 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A2 = CLBLM_R_X13Y102_SLICE_X19Y102_DO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A4 = CLBLM_R_X15Y100_SLICE_X20Y100_DO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A5 = CLBLM_R_X15Y101_SLICE_X20Y101_AO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_A6 = CLBLM_R_X15Y100_SLICE_X20Y100_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B1 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B5 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_B6 = 1'b1;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C2 = CLBLM_R_X15Y100_SLICE_X21Y100_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D1 = 1'b1;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D2 = CLBLM_R_X15Y101_SLICE_X20Y101_BO5;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C4 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = 1'b1;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C5 = CLBLM_L_X16Y108_SLICE_X22Y108_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_D4 = CLBLM_R_X15Y102_SLICE_X20Y102_CO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_C6 = CLBLM_L_X16Y102_SLICE_X23Y102_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y100_SLICE_X20Y100_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D1 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D2 = CLBLM_L_X16Y102_SLICE_X22Y102_BO5;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D3 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D4 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D5 = 1'b1;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_D6 = CLBLM_R_X15Y103_SLICE_X20Y103_DO6;
  assign CLBLM_L_X16Y104_SLICE_X22Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLM_R_X15Y115_SLICE_X20Y115_AQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLM_R_X15Y116_SLICE_X20Y116_BQ;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A1 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A2 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A3 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A4 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B1 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B2 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B3 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B4 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_B6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C1 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C2 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C4 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C5 = CLBLM_R_X15Y101_SLICE_X21Y101_AO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_C6 = CLBLM_R_X13Y101_SLICE_X19Y101_BO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D1 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D2 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D4 = CLBLM_R_X13Y101_SLICE_X19Y101_CO6;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y101_SLICE_X21Y101_D6 = CLBLM_R_X15Y101_SLICE_X21Y101_BO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A1 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A2 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A5 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_A6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B1 = CLBLM_R_X13Y101_SLICE_X19Y101_DO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B2 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B3 = CLBLM_R_X13Y100_SLICE_X18Y100_CO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B5 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_B6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C1 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C2 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C3 = CLBLM_L_X12Y101_SLICE_X17Y101_BO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C4 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C5 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_C6 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_D = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_D = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C5 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C6 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D1 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D2 = 1'b1;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D3 = CLBLM_R_X15Y101_SLICE_X21Y101_BO5;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X15Y101_SLICE_X20Y101_D6 = CLBLM_R_X15Y101_SLICE_X20Y101_BO6;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A2 = CLBLM_L_X12Y103_SLICE_X17Y103_BO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A5 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_A6 = 1'b1;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B1 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B2 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B3 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B4 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B5 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_B6 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C5 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_C6 = CLBLM_L_X12Y103_SLICE_X17Y103_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D1 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D2 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A4 = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D4 = CLBLM_R_X15Y102_SLICE_X21Y102_AO5;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D5 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X15Y102_SLICE_X21Y102_D6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A5 = CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A6 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A1 = CLBLM_R_X15Y102_SLICE_X20Y102_DO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A3 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A4 = CLBLM_R_X15Y103_SLICE_X20Y103_BO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A5 = 1'b1;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_A6 = CLBLM_R_X15Y101_SLICE_X20Y101_DO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B2 = CLBLM_R_X13Y101_SLICE_X19Y101_AO5;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B3 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B5 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_B6 = CLBLM_L_X12Y103_SLICE_X17Y103_CO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C2 = CLBLM_L_X12Y103_SLICE_X17Y103_CO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C3 = CLBLM_R_X13Y101_SLICE_X19Y101_AO5;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C4 = 1'b1;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C5 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_C6 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_D = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D1 = 1'b1;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D2 = CLBLM_R_X15Y101_SLICE_X21Y101_AO5;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D3 = 1'b1;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_D6 = CLBLM_R_X15Y102_SLICE_X20Y102_BO6;
  assign CLBLM_R_X15Y102_SLICE_X20Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C2 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = 1'b0;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A1 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A3 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A4 = CLBLM_R_X15Y102_SLICE_X21Y102_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_A6 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B1 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B3 = CLBLM_R_X15Y103_SLICE_X20Y103_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B4 = CLBLM_L_X16Y110_SLICE_X23Y110_DO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_B6 = CLBLM_R_X15Y103_SLICE_X21Y103_AO5;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C1 = CLBLM_R_X15Y102_SLICE_X21Y102_CO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C2 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C4 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C5 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_C6 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLM_L_X16Y115_SLICE_X22Y115_AQ;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D1 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D2 = CLBLM_R_X15Y103_SLICE_X20Y103_AO5;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D3 = CLBLM_R_X15Y103_SLICE_X20Y103_DO6;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D4 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D5 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X21Y103_D6 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A1 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A2 = CLBLM_R_X13Y100_SLICE_X19Y100_AO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A3 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A4 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A5 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_A6 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLM_R_X15Y115_SLICE_X21Y115_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B1 = CLBLM_R_X15Y102_SLICE_X21Y102_DO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B5 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_B6 = CLBLM_R_X13Y102_SLICE_X19Y102_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C4 = CLBLM_L_X12Y101_SLICE_X17Y101_AO6;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C5 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_C6 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D1 = CLBLM_R_X15Y102_SLICE_X20Y102_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D2 = CLBLM_R_X13Y103_SLICE_X19Y103_AO5;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D3 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D4 = CLBLM_L_X12Y101_SLICE_X17Y101_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D5 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_R_X15Y103_SLICE_X20Y103_D6 = CLBLM_R_X15Y100_SLICE_X20Y100_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A1 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A2 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A3 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A4 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A5 = CLBLM_R_X11Y102_SLICE_X14Y102_BO6;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_A6 = CLBLM_L_X12Y102_SLICE_X17Y102_AO5;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_B6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_C6 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X17Y100_D6 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_A6 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_C6 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D1 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D2 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D3 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D4 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D5 = 1'b1;
  assign CLBLM_L_X12Y100_SLICE_X16Y100_D6 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A1 = CLBLM_R_X15Y103_SLICE_X21Y103_DO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A2 = CLBLM_L_X16Y104_SLICE_X22Y104_CO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A3 = CLBLM_R_X15Y103_SLICE_X21Y103_AO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A4 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A5 = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B2 = CLBLM_R_X15Y100_SLICE_X21Y100_BO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B4 = CLBLM_R_X15Y103_SLICE_X21Y103_AO5;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B5 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_B6 = CLBLM_R_X15Y104_SLICE_X21Y104_CO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C2 = CLBLM_R_X15Y103_SLICE_X20Y103_CO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C3 = CLBLM_R_X15Y108_SLICE_X21Y108_CO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C4 = CLBLM_L_X16Y110_SLICE_X23Y110_DO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D1 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D2 = CLBLM_L_X16Y103_SLICE_X22Y103_CO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D3 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D4 = CLBLM_R_X15Y109_SLICE_X21Y109_BO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D5 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X15Y104_SLICE_X21Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A2 = CLBLM_R_X15Y102_SLICE_X20Y102_BO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A3 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A4 = CLBLM_R_X15Y104_SLICE_X20Y104_BO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_A6 = CLBLM_R_X15Y102_SLICE_X21Y102_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B1 = CLBLM_R_X15Y108_SLICE_X20Y108_DO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B5 = CLBLM_R_X13Y102_SLICE_X19Y102_BO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_B6 = CLBLM_R_X15Y109_SLICE_X20Y109_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C4 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C5 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_C6 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D1 = CLBLM_L_X16Y103_SLICE_X23Y103_AO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D2 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D4 = CLBLM_R_X15Y101_SLICE_X20Y101_CO6;
  assign CLBLM_R_X15Y104_SLICE_X20Y104_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A1 = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A2 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A3 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A4 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A5 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_A6 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B1 = CLBLM_R_X13Y100_SLICE_X18Y100_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B2 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B3 = CLBLM_L_X12Y101_SLICE_X16Y101_AO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B4 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B5 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_B6 = CLBLM_R_X11Y101_SLICE_X14Y101_BO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C1 = CLBLM_R_X13Y102_SLICE_X18Y102_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C2 = CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C3 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C5 = CLBLM_L_X12Y101_SLICE_X17Y101_DO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_C6 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D2 = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D3 = CLBLM_R_X11Y101_SLICE_X15Y101_AO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D4 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D5 = 1'b1;
  assign CLBLM_L_X12Y101_SLICE_X17Y101_D6 = 1'b1;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A1 = CLBLM_L_X10Y100_SLICE_X12Y100_BO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A3 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A4 = CLBLM_R_X11Y100_SLICE_X14Y100_BO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A5 = 1'b1;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_A6 = 1'b1;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B1 = CLBLM_L_X12Y101_SLICE_X16Y101_DO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B4 = 1'b1;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B5 = CLBLM_R_X11Y102_SLICE_X15Y102_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_B6 = CLBLM_L_X12Y101_SLICE_X16Y101_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C1 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C2 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C3 = CLBLM_L_X12Y103_SLICE_X16Y103_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C4 = CLBLM_L_X12Y101_SLICE_X16Y101_AO5;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C5 = CLBLM_R_X11Y101_SLICE_X15Y101_AO5;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D1 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D2 = 1'b1;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D3 = CLBLM_R_X11Y101_SLICE_X14Y101_DO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D5 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X12Y101_SLICE_X16Y101_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A1 = CLBLM_R_X15Y105_SLICE_X21Y105_DO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A2 = CLBLM_L_X16Y105_SLICE_X22Y105_CO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A3 = CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A5 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_A6 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B1 = CLBLM_L_X16Y103_SLICE_X23Y103_CO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B2 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B3 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B4 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B5 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_B6 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C1 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C2 = CLBLM_R_X15Y102_SLICE_X21Y102_BO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C5 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_C6 = CLBLM_R_X15Y104_SLICE_X20Y104_CO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D1 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D2 = CLBLM_L_X16Y104_SLICE_X23Y104_CO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D4 = CLBLM_R_X15Y105_SLICE_X21Y105_CO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B3 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D5 = CLBLM_R_X15Y105_SLICE_X21Y105_BO5;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_D6 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B4 = CLBLM_L_X16Y110_SLICE_X22Y110_DO6;
  assign CLBLM_R_X15Y105_SLICE_X21Y105_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A1 = CLBLM_L_X16Y101_SLICE_X22Y101_AQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B5 = CLBLM_L_X16Y105_SLICE_X23Y105_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A2 = CLBLM_R_X15Y102_SLICE_X21Y102_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A4 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_A6 = CLBLM_L_X16Y102_SLICE_X22Y102_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = 1'b1;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B1 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B2 = CLBLM_R_X15Y101_SLICE_X20Y101_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B5 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_B6 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C4 = CLBLM_R_X15Y102_SLICE_X21Y102_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_C5 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D1 = CLBLM_R_X15Y105_SLICE_X21Y105_BO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D3 = CLBLM_L_X16Y103_SLICE_X22Y103_CO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C2 = CLBLM_L_X16Y105_SLICE_X23Y105_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_R_X15Y105_SLICE_X20Y105_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C4 = CLBLM_L_X16Y110_SLICE_X22Y110_DO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C5 = CLBLM_L_X16Y105_SLICE_X22Y105_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_C6 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLM_L_X16Y115_SLICE_X23Y115_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_L_X16Y115_SLICE_X23Y115_AQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D2 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D3 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D5 = CLBLM_R_X15Y105_SLICE_X20Y105_CO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A1 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A2 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A3 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_A6 = 1'b1;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_D6 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B1 = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B2 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B3 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_B6 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C2 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C3 = CLBLM_R_X11Y102_SLICE_X14Y102_AO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C4 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C5 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_C6 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X16Y105_SLICE_X22Y105_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D2 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D3 = CLBLM_R_X11Y102_SLICE_X14Y102_AO6;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D4 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D5 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y102_SLICE_X17Y102_D6 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A1 = CLBLM_L_X12Y102_SLICE_X16Y102_DO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A2 = CLBLM_R_X11Y102_SLICE_X14Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A3 = CLBLM_R_X11Y101_SLICE_X14Y101_AQ;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A5 = CLBLM_R_X11Y103_SLICE_X15Y103_AO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B1 = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B2 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B3 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B4 = CLBLM_R_X11Y101_SLICE_X15Y101_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_CO5;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y132_SLICE_X21Y132_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C2 = CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C4 = CLBLM_L_X12Y102_SLICE_X16Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C5 = CLBLM_R_X11Y102_SLICE_X15Y102_AO5;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_C6 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D1 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D2 = CLBLM_R_X11Y100_SLICE_X14Y100_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D3 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D4 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D5 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_D6 = 1'b1;
  assign CLBLM_L_X12Y102_SLICE_X16Y102_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_A6 = 1'b1;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A1 = CLBLM_R_X15Y105_SLICE_X20Y105_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A2 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A4 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A5 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_A6 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B1 = CLBLM_R_X15Y101_SLICE_X21Y101_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B2 = CLBLM_L_X16Y105_SLICE_X23Y105_AO5;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B3 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B4 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B5 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = 1'b1;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_B6 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C1 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C2 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C3 = CLBLM_R_X15Y101_SLICE_X21Y101_DO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C4 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C5 = CLBLM_R_X15Y105_SLICE_X21Y105_AO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_C6 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D1 = CLBLM_R_X15Y106_SLICE_X21Y106_AO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D4 = CLBLM_R_X15Y106_SLICE_X21Y106_CO6;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D5 = 1'b1;
  assign CLBLM_R_X15Y106_SLICE_X21Y106_D6 = CLBLM_R_X15Y112_SLICE_X21Y112_CO5;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A3 = CLBLM_R_X15Y105_SLICE_X20Y105_AO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A4 = CLBLM_R_X15Y106_SLICE_X20Y106_BO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A5 = CLBLM_L_X16Y105_SLICE_X23Y105_AO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_A6 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B1 = CLBLM_R_X15Y104_SLICE_X20Y104_DO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B3 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B4 = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B5 = CLBLM_R_X15Y109_SLICE_X20Y109_CO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C1 = 1'b1;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C1 = CLBLM_R_X15Y105_SLICE_X20Y105_AO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C3 = CLBLM_R_X15Y104_SLICE_X20Y104_DO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_C6 = CLBLM_R_X15Y109_SLICE_X20Y109_BO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C2 = 1'b1;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D1 = CLBLM_R_X15Y100_SLICE_X21Y100_AO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D3 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D5 = CLBLM_L_X16Y104_SLICE_X23Y104_AQ;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_D6 = CLBLM_L_X16Y109_SLICE_X23Y109_BO6;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C5 = 1'b1;
  assign CLBLM_R_X15Y132_SLICE_X20Y132_C6 = 1'b1;
  assign CLBLM_R_X15Y106_SLICE_X20Y106_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A2 = CLBLM_L_X16Y126_SLICE_X23Y126_BO5;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_A4 = CLBLM_R_X13Y124_SLICE_X18Y124_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A1 = CLBLM_L_X12Y103_SLICE_X17Y103_DO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A2 = CLBLM_R_X13Y103_SLICE_X18Y103_CO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A3 = CLBLM_L_X12Y102_SLICE_X17Y102_BO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A5 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_A6 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B2 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B3 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B4 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_B6 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C2 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C3 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C4 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C5 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_C6 = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D1 = 1'b1;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D2 = CLBLM_R_X13Y101_SLICE_X18Y101_AQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D3 = CLBLM_L_X12Y103_SLICE_X16Y103_DO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_D6 = 1'b1;
  assign CLBLM_L_X12Y103_SLICE_X17Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A1 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A2 = CLBLM_R_X11Y103_SLICE_X15Y103_CO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A3 = CLBLM_L_X12Y102_SLICE_X16Y102_DO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A4 = CLBLM_L_X12Y103_SLICE_X16Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_A6 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B2 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B4 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B5 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_B6 = 1'b1;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C4 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_C6 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D1 = CLBLM_L_X12Y102_SLICE_X16Y102_AQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D2 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D4 = CLBLM_L_X12Y101_SLICE_X16Y101_BQ;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D5 = 1'b1;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_D6 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X12Y103_SLICE_X16Y103_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_C5 = CLBLM_L_X16Y126_SLICE_X22Y126_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = CLBLM_L_X16Y126_SLICE_X23Y126_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A1 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A2 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A3 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A4 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A5 = CLBLM_R_X15Y105_SLICE_X20Y105_CO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_A6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B1 = CLBLM_R_X15Y107_SLICE_X21Y107_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B2 = CLBLM_R_X15Y107_SLICE_X20Y107_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B4 = CLBLM_R_X15Y108_SLICE_X21Y108_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B5 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C1 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C2 = CLBLM_R_X15Y107_SLICE_X20Y107_CO5;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C3 = CLBLM_R_X15Y106_SLICE_X21Y106_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C5 = CLBLM_R_X15Y108_SLICE_X21Y108_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_C6 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D1 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D3 = CLBLM_L_X16Y107_SLICE_X23Y107_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D4 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D5 = CLBLM_R_X15Y107_SLICE_X21Y107_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_D6 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X15Y107_SLICE_X21Y107_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A1 = CLBLM_R_X15Y107_SLICE_X20Y107_BO5;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A3 = CLBLM_R_X15Y107_SLICE_X20Y107_DO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A4 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A5 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A5 = CLBLM_L_X16Y107_SLICE_X23Y107_AO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_A6 = CLBLM_R_X15Y107_SLICE_X20Y107_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A6 = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B1 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B2 = CLBLM_R_X15Y105_SLICE_X20Y105_BO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B3 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B4 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B5 = CLBLM_L_X16Y106_SLICE_X22Y106_BO5;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_B6 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C1 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C2 = CLBLM_R_X15Y107_SLICE_X21Y107_AO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X16Y126_SLICE_X22Y126_D6 = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C4 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_C6 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D1 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D2 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D3 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D4 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D5 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = 1'b1;
  assign CLBLM_R_X15Y107_SLICE_X20Y107_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A3 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A4 = CLBLM_L_X12Y103_SLICE_X16Y103_BO5;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A5 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A6 = CLBLM_L_X12Y102_SLICE_X16Y102_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B1 = CLBLM_R_X11Y101_SLICE_X14Y101_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B2 = CLBLM_L_X12Y103_SLICE_X16Y103_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B3 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B4 = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C1 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C2 = CLBLM_L_X12Y101_SLICE_X17Y101_DO5;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C3 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C5 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C6 = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D1 = CLBLM_L_X12Y102_SLICE_X16Y102_BQ;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D4 = CLBLM_L_X12Y103_SLICE_X16Y103_BO5;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D5 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D6 = CLBLM_L_X12Y101_SLICE_X17Y101_DO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_L_X16Y114_SLICE_X23Y114_AQ;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A5 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B1 = CLBLM_R_X15Y107_SLICE_X21Y107_CQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B2 = CLBLM_R_X15Y106_SLICE_X21Y106_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B4 = CLBLM_R_X15Y112_SLICE_X21Y112_DO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_B6 = CLBLM_R_X15Y109_SLICE_X21Y109_CO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C2 = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C3 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C4 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D1 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D2 = 1'b1;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D3 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D4 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D5 = CLBLM_R_X15Y109_SLICE_X21Y109_DO6;
  assign CLBLM_R_X15Y108_SLICE_X21Y108_D6 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A1 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A2 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A3 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A4 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A5 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_A6 = 1'b1;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B5 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C4 = 1'b1;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_C6 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D1 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D2 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D4 = CLBLM_R_X15Y108_SLICE_X20Y108_AO5;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D5 = 1'b1;
  assign CLBLM_R_X15Y108_SLICE_X20Y108_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A2 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A3 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A4 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A5 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_A6 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B2 = CLBLM_L_X16Y109_SLICE_X23Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B4 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B5 = CLBLM_R_X15Y109_SLICE_X21Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_B6 = CLBLM_L_X16Y109_SLICE_X23Y109_BO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C1 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C2 = CLBLM_R_X15Y107_SLICE_X21Y107_CQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C3 = CLBLM_L_X16Y109_SLICE_X22Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C4 = CLBLM_L_X16Y109_SLICE_X22Y109_DO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D1 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D3 = CLBLM_L_X16Y109_SLICE_X22Y109_AO6;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D4 = CLBLM_L_X16Y109_SLICE_X23Y109_AO5;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X21Y109_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A3 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B1 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C2 = CLBLM_R_X15Y109_SLICE_X21Y109_AO5;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C4 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C5 = CLBLM_L_X16Y109_SLICE_X22Y109_CO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D1 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D2 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D3 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D4 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D5 = 1'b1;
  assign CLBLM_R_X15Y109_SLICE_X20Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A1 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A2 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A3 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A4 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A5 = CLBLM_L_X12Y103_SLICE_X17Y103_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A1 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A2 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A3 = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A4 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A5 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B1 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B3 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B4 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B5 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B6 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C1 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C2 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C3 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C4 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C5 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C6 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D3 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D4 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D6 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A2 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A3 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A4 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A5 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_A6 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B2 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B3 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B4 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B5 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_B6 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C1 = CLBLM_L_X16Y109_SLICE_X22Y109_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C3 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C4 = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_C6 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D1 = CLBLM_R_X15Y110_SLICE_X21Y110_AO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D2 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D3 = CLBLM_R_X15Y106_SLICE_X20Y106_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D4 = CLBLM_R_X15Y110_SLICE_X20Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D5 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X21Y110_D6 = CLBLM_L_X16Y105_SLICE_X22Y105_AQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B3 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A2 = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A3 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A4 = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_B4 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_A6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_R_X15Y116_SLICE_X21Y116_AQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B2 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B3 = CLBLM_R_X15Y104_SLICE_X21Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B4 = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B5 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_B6 = CLBLM_R_X13Y104_SLICE_X19Y104_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C1 = CLBLM_R_X15Y104_SLICE_X20Y104_AQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C4 = CLBLM_R_X15Y108_SLICE_X20Y108_AO5;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_C6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_R_X15Y114_SLICE_X20Y114_AQ;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D1 = 1'b1;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D4 = CLBLM_L_X16Y109_SLICE_X23Y109_AO5;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X15Y110_SLICE_X20Y110_D6 = CLBLM_R_X15Y107_SLICE_X21Y107_BQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C2 = CLBLM_R_X15Y107_SLICE_X20Y107_AQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C3 = CLBLM_L_X16Y106_SLICE_X23Y106_BO5;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_C6 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A2 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A4 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A6 = 1'b1;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D4 = CLBLM_L_X16Y104_SLICE_X22Y104_BQ;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D5 = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B6 = 1'b1;
  assign CLBLM_L_X16Y106_SLICE_X22Y106_D6 = CLBLM_L_X16Y108_SLICE_X22Y108_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A4 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A1 = CLBLM_R_X15Y112_SLICE_X20Y112_DO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A3 = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A4 = CLBLM_R_X15Y111_SLICE_X21Y111_BO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A5 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_A6 = CLBLM_R_X15Y111_SLICE_X21Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B1 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B3 = CLBLM_R_X15Y111_SLICE_X20Y111_AO5;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B4 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B5 = CLBLM_R_X15Y110_SLICE_X21Y110_CO5;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_B6 = CLBLM_L_X16Y109_SLICE_X23Y109_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C1 = CLBLM_L_X16Y104_SLICE_X22Y104_AQ;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C2 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C3 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C4 = CLBLM_L_X16Y109_SLICE_X23Y109_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C5 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D1 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D4 = CLBLM_R_X15Y110_SLICE_X20Y110_AO5;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D5 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_D6 = CLBLM_R_X15Y110_SLICE_X21Y110_AO5;
  assign CLBLM_R_X15Y111_SLICE_X21Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A1 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A2 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A4 = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A5 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_A6 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B1 = CLBLM_L_X12Y116_SLICE_X17Y116_AQ;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B3 = CLBLM_R_X15Y111_SLICE_X21Y111_DO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B4 = CLBLM_R_X13Y114_SLICE_X18Y114_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_B6 = CLBLM_R_X15Y111_SLICE_X20Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C1 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C2 = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C3 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C4 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C5 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_C6 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D1 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D2 = CLBLM_R_X15Y110_SLICE_X21Y110_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D3 = 1'b1;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D4 = CLBLM_L_X12Y116_SLICE_X17Y116_A5Q;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D5 = CLBLM_R_X13Y115_SLICE_X18Y115_CO6;
  assign CLBLM_R_X15Y111_SLICE_X20Y111_D6 = CLBLM_R_X13Y111_SLICE_X19Y111_BO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A2 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A3 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A4 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B1 = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B3 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B4 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B5 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B6 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_A5Q;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C1 = CLBLM_L_X12Y104_SLICE_X16Y104_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C3 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C6 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D1 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D2 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D5 = CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A1 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A2 = CLBLM_L_X10Y104_SLICE_X13Y104_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A3 = CLBLM_R_X11Y104_SLICE_X14Y104_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A4 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A5 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B1 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B2 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B5 = CLBLM_L_X12Y104_SLICE_X16Y104_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C1 = CLBLM_R_X11Y103_SLICE_X14Y103_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A2 = CLBLM_R_X15Y110_SLICE_X21Y110_BO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A4 = CLBLM_R_X15Y112_SLICE_X21Y112_BO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A5 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_A6 = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B1 = CLBLM_R_X15Y104_SLICE_X21Y104_BQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_B6 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C1 = CLBLM_L_X16Y106_SLICE_X22Y106_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C4 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C5 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_C6 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D1 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D4 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_D6 = CLBLM_L_X8Y111_SLICE_X10Y111_BQ;
  assign CLBLM_R_X15Y112_SLICE_X21Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A1 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A2 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A3 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A4 = CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A5 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_A6 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B1 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B2 = CLBLM_L_X16Y111_SLICE_X22Y111_BQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B3 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B4 = CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_B6 = CLBLM_L_X12Y115_SLICE_X17Y115_A5Q;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A6 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C1 = CLBLM_R_X15Y112_SLICE_X20Y112_AO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C2 = CLBLM_L_X16Y111_SLICE_X22Y111_AQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C3 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C4 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C5 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_C6 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D1 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D2 = CLBLM_R_X15Y111_SLICE_X21Y111_AQ;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D3 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D4 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D5 = 1'b1;
  assign CLBLM_R_X15Y112_SLICE_X20Y112_D6 = CLBLM_R_X15Y113_SLICE_X20Y113_AO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C1 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C2 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C3 = CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_R_X15Y117_SLICE_X21Y117_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C5 = CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A1 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A3 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A4 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A6 = CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_L_X16Y117_SLICE_X22Y117_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B1 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B3 = CLBLM_L_X12Y103_SLICE_X16Y103_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B4 = CLBLM_R_X15Y112_SLICE_X21Y112_BO5;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B5 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B6 = CLBLM_L_X16Y110_SLICE_X23Y110_AO5;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C4 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C5 = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D1 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D2 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A1 = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A2 = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A3 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B4 = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C1 = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C2 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C3 = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C4 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C6 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D1 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D2 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D3 = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D4 = CLBLM_L_X12Y111_SLICE_X16Y111_AO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D5 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D6 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A2 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A3 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A4 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A5 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_A6 = CLBLM_R_X15Y115_SLICE_X21Y115_BO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B3 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B4 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B5 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_B6 = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C1 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C2 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C3 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C4 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C5 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_C6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D1 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D2 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D3 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D4 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D5 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X21Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A1 = CLBLM_R_X13Y111_SLICE_X18Y111_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A2 = CLBLM_L_X16Y110_SLICE_X22Y110_AQ;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A3 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A4 = CLBLM_L_X16Y111_SLICE_X23Y111_AQ;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A5 = CLBLM_R_X15Y112_SLICE_X21Y112_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_A6 = CLBLM_R_X13Y111_SLICE_X18Y111_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B1 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B2 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B3 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B4 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B5 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_B6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C1 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C2 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C3 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C4 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C5 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_C6 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D1 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D2 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D3 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D4 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D5 = 1'b1;
  assign CLBLM_R_X15Y113_SLICE_X20Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y115_SLICE_X3Y115_A5Q;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X15Y105_SLICE_X21Y105_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = CLBLM_R_X3Y115_SLICE_X2Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = CLBLM_R_X13Y111_SLICE_X19Y111_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A1 = CLBLM_R_X15Y114_SLICE_X21Y114_DO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A2 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_A6 = CLBLM_R_X15Y112_SLICE_X21Y112_CO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B1 = CLBLM_R_X15Y115_SLICE_X21Y115_BO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B2 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B4 = CLBLM_R_X11Y110_SLICE_X14Y110_BQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B5 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_B6 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C1 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C3 = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_C6 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D2 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D5 = CLBLM_L_X16Y113_SLICE_X22Y113_BO5;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_D6 = CLBLM_R_X15Y114_SLICE_X21Y114_AQ;
  assign CLBLM_R_X15Y114_SLICE_X21Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A1 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A2 = CLBLM_R_X15Y114_SLICE_X21Y114_BO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A4 = CLBLM_L_X16Y114_SLICE_X23Y114_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A5 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_A6 = CLBLM_R_X15Y114_SLICE_X20Y114_CO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B1 = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B2 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B4 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_B6 = 1'b1;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C2 = CLBLM_R_X15Y114_SLICE_X20Y114_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_C6 = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D1 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D2 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D4 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X15Y114_SLICE_X20Y114_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A2 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A4 = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A5 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A6 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B1 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B5 = CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B6 = CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C1 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C4 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C5 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C6 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D1 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D3 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D5 = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D6 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A1 = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A2 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A4 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A5 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A6 = 1'b1;
  assign CLBLM_R_X13Y123_SLICE_X19Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B1 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B3 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C1 = CLBLM_L_X12Y111_SLICE_X17Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C5 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C6 = CLBLM_L_X12Y110_SLICE_X16Y110_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D4 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D5 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_L_X16Y118_SLICE_X23Y118_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A1 = CLBLM_R_X15Y115_SLICE_X20Y115_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A2 = CLBLM_R_X15Y115_SLICE_X20Y115_BO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A5 = CLBLM_R_X15Y115_SLICE_X21Y115_CO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_A6 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B2 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B4 = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_B6 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C1 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C2 = CLBLM_R_X15Y115_SLICE_X21Y115_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C5 = CLBLM_R_X15Y114_SLICE_X21Y114_CO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_C6 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D2 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D4 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D5 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_D6 = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_R_X15Y115_SLICE_X21Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A1 = CLBLM_R_X15Y115_SLICE_X20Y115_BO5;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A4 = CLBLM_R_X15Y116_SLICE_X20Y116_BQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A5 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_A6 = CLBLM_R_X15Y115_SLICE_X20Y115_CO6;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B3 = CLBLM_L_X16Y107_SLICE_X22Y107_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B1 = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B2 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B4 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_B6 = 1'b1;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C1 = CLBLM_R_X15Y114_SLICE_X20Y114_BO6;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C2 = CLBLM_R_X15Y115_SLICE_X20Y115_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_C6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D1 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D2 = CLBLM_R_X15Y116_SLICE_X20Y116_BQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D4 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_D6 = CLBLM_R_X15Y114_SLICE_X20Y114_BO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLM_R_X15Y115_SLICE_X20Y115_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C1 = CLBLM_L_X16Y107_SLICE_X23Y107_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = 1'b1;
  assign CLBLM_L_X16Y107_SLICE_X22Y107_C3 = CLBLM_L_X16Y106_SLICE_X23Y106_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A1 = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A2 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A4 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A5 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A6 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B1 = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B2 = CLBLM_R_X11Y114_SLICE_X15Y114_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B4 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B5 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B6 = CLBLM_R_X11Y114_SLICE_X14Y114_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C1 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C2 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C3 = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C4 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C6 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D1 = CLBLM_R_X13Y111_SLICE_X18Y111_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D4 = CLBLM_L_X12Y111_SLICE_X17Y111_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D5 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D6 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A1 = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A2 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A3 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A6 = CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B1 = CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B2 = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B3 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B4 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B6 = CLBLM_R_X11Y117_SLICE_X15Y117_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C1 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C2 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C4 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C5 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C6 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D2 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D3 = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D5 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A1 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A4 = CLBLM_R_X15Y113_SLICE_X21Y113_AO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A5 = CLBLM_R_X15Y114_SLICE_X20Y114_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_A6 = CLBLM_R_X15Y116_SLICE_X21Y116_CO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B1 = CLBLM_R_X15Y116_SLICE_X21Y116_DO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B3 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B4 = CLBLM_R_X15Y116_SLICE_X21Y116_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_B6 = CLBLM_R_X13Y114_SLICE_X19Y114_AO5;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C1 = CLBLM_L_X16Y116_SLICE_X23Y116_DO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C2 = CLBLM_R_X15Y116_SLICE_X21Y116_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C4 = CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C5 = CLBLM_R_X13Y114_SLICE_X19Y114_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_C6 = CLBLM_R_X15Y113_SLICE_X21Y113_BO6;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D1 = CLBLM_R_X15Y116_SLICE_X21Y116_BQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D3 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D4 = CLBLM_L_X16Y116_SLICE_X22Y116_BO5;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_D6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y116_SLICE_X21Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A1 = CLBLM_R_X15Y116_SLICE_X20Y116_DO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A3 = CLBLM_L_X16Y116_SLICE_X23Y116_BQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A4 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_A6 = CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B1 = CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B3 = CLBLM_R_X15Y116_SLICE_X20Y116_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B4 = CLBLM_R_X15Y115_SLICE_X20Y115_DO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_B6 = CLBLM_R_X15Y116_SLICE_X20Y116_CO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C2 = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C3 = CLBLM_R_X15Y114_SLICE_X20Y114_DO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C4 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C5 = 1'b1;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_C6 = 1'b1;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D1 = CLBLM_R_X15Y116_SLICE_X20Y116_CO5;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D2 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D5 = CLBLM_R_X15Y131_SLICE_X20Y131_B5Q;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_D6 = CLBLM_R_X15Y116_SLICE_X20Y116_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X15Y116_SLICE_X20Y116_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = 1'b1;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_O = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A1 = CLBLM_R_X11Y112_SLICE_X14Y112_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A2 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_SR = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A4 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B1 = CLBLM_L_X12Y113_SLICE_X16Y113_A5Q;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B2 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B4 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B5 = CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C3 = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_A5Q;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D1 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A1 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A2 = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A3 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A4 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A5 = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B1 = CLBLM_R_X11Y113_SLICE_X15Y113_A5Q;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B3 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B4 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B5 = CLBLM_L_X10Y117_SLICE_X13Y117_A5Q;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C1 = CLBLM_R_X13Y120_SLICE_X18Y120_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C3 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C4 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C6 = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D1 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D2 = CLBLM_L_X12Y113_SLICE_X17Y113_AO5;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D3 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
endmodule
