module top(
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  input RIOB33_X105Y77_IOB_X1Y78_IPAD,
  output LIOB33_SING_X0Y0_IOB_X0Y0_OPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_SING_X0Y200_IOB_X0Y200_OPAD,
  output LIOB33_SING_X0Y249_IOB_X0Y249_OPAD,
  output LIOB33_SING_X0Y50_IOB_X0Y50_OPAD,
  output LIOB33_SING_X0Y99_IOB_X0Y99_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y1_IOB_X0Y1_OPAD,
  output LIOB33_X0Y1_IOB_X0Y2_OPAD,
  output LIOB33_X0Y201_IOB_X0Y201_OPAD,
  output LIOB33_X0Y201_IOB_X0Y202_OPAD,
  output LIOB33_X0Y203_IOB_X0Y203_OPAD,
  output LIOB33_X0Y203_IOB_X0Y204_OPAD,
  output LIOB33_X0Y205_IOB_X0Y205_OPAD,
  output LIOB33_X0Y205_IOB_X0Y206_OPAD,
  output LIOB33_X0Y207_IOB_X0Y207_OPAD,
  output LIOB33_X0Y207_IOB_X0Y208_OPAD,
  output LIOB33_X0Y209_IOB_X0Y209_OPAD,
  output LIOB33_X0Y209_IOB_X0Y210_OPAD,
  output LIOB33_X0Y211_IOB_X0Y211_OPAD,
  output LIOB33_X0Y211_IOB_X0Y212_OPAD,
  output LIOB33_X0Y213_IOB_X0Y213_OPAD,
  output LIOB33_X0Y213_IOB_X0Y214_OPAD,
  output LIOB33_X0Y215_IOB_X0Y215_OPAD,
  output LIOB33_X0Y215_IOB_X0Y216_OPAD,
  output LIOB33_X0Y217_IOB_X0Y217_OPAD,
  output LIOB33_X0Y217_IOB_X0Y218_OPAD,
  output LIOB33_X0Y219_IOB_X0Y219_OPAD,
  output LIOB33_X0Y219_IOB_X0Y220_OPAD,
  output LIOB33_X0Y221_IOB_X0Y221_OPAD,
  output LIOB33_X0Y221_IOB_X0Y222_OPAD,
  output LIOB33_X0Y223_IOB_X0Y223_OPAD,
  output LIOB33_X0Y223_IOB_X0Y224_OPAD,
  output LIOB33_X0Y225_IOB_X0Y225_OPAD,
  output LIOB33_X0Y225_IOB_X0Y226_OPAD,
  output LIOB33_X0Y227_IOB_X0Y227_OPAD,
  output LIOB33_X0Y227_IOB_X0Y228_OPAD,
  output LIOB33_X0Y229_IOB_X0Y229_OPAD,
  output LIOB33_X0Y229_IOB_X0Y230_OPAD,
  output LIOB33_X0Y231_IOB_X0Y231_OPAD,
  output LIOB33_X0Y231_IOB_X0Y232_OPAD,
  output LIOB33_X0Y233_IOB_X0Y233_OPAD,
  output LIOB33_X0Y233_IOB_X0Y234_OPAD,
  output LIOB33_X0Y235_IOB_X0Y235_OPAD,
  output LIOB33_X0Y235_IOB_X0Y236_OPAD,
  output LIOB33_X0Y237_IOB_X0Y237_OPAD,
  output LIOB33_X0Y237_IOB_X0Y238_OPAD,
  output LIOB33_X0Y239_IOB_X0Y239_OPAD,
  output LIOB33_X0Y239_IOB_X0Y240_OPAD,
  output LIOB33_X0Y241_IOB_X0Y241_OPAD,
  output LIOB33_X0Y241_IOB_X0Y242_OPAD,
  output LIOB33_X0Y243_IOB_X0Y243_OPAD,
  output LIOB33_X0Y243_IOB_X0Y244_OPAD,
  output LIOB33_X0Y245_IOB_X0Y245_OPAD,
  output LIOB33_X0Y245_IOB_X0Y246_OPAD,
  output LIOB33_X0Y247_IOB_X0Y247_OPAD,
  output LIOB33_X0Y247_IOB_X0Y248_OPAD,
  output LIOB33_X0Y3_IOB_X0Y3_OPAD,
  output LIOB33_X0Y3_IOB_X0Y4_OPAD,
  output LIOB33_X0Y51_IOB_X0Y51_OPAD,
  output LIOB33_X0Y51_IOB_X0Y52_OPAD,
  output LIOB33_X0Y53_IOB_X0Y53_OPAD,
  output LIOB33_X0Y53_IOB_X0Y54_OPAD,
  output LIOB33_X0Y55_IOB_X0Y55_OPAD,
  output LIOB33_X0Y55_IOB_X0Y56_OPAD,
  output LIOB33_X0Y57_IOB_X0Y57_OPAD,
  output LIOB33_X0Y57_IOB_X0Y58_OPAD,
  output LIOB33_X0Y59_IOB_X0Y59_OPAD,
  output LIOB33_X0Y59_IOB_X0Y60_OPAD,
  output LIOB33_X0Y5_IOB_X0Y5_OPAD,
  output LIOB33_X0Y5_IOB_X0Y6_OPAD,
  output LIOB33_X0Y61_IOB_X0Y61_OPAD,
  output LIOB33_X0Y61_IOB_X0Y62_OPAD,
  output LIOB33_X0Y63_IOB_X0Y63_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output LIOB33_X0Y67_IOB_X0Y67_OPAD,
  output LIOB33_X0Y67_IOB_X0Y68_OPAD,
  output LIOB33_X0Y69_IOB_X0Y69_OPAD,
  output LIOB33_X0Y69_IOB_X0Y70_OPAD,
  output LIOB33_X0Y71_IOB_X0Y71_OPAD,
  output LIOB33_X0Y71_IOB_X0Y72_OPAD,
  output LIOB33_X0Y73_IOB_X0Y73_OPAD,
  output LIOB33_X0Y73_IOB_X0Y74_OPAD,
  output LIOB33_X0Y75_IOB_X0Y75_OPAD,
  output LIOB33_X0Y75_IOB_X0Y76_OPAD,
  output LIOB33_X0Y77_IOB_X0Y77_OPAD,
  output LIOB33_X0Y77_IOB_X0Y78_OPAD,
  output LIOB33_X0Y79_IOB_X0Y79_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output LIOB33_X0Y81_IOB_X0Y81_OPAD,
  output LIOB33_X0Y81_IOB_X0Y82_OPAD,
  output LIOB33_X0Y83_IOB_X0Y83_OPAD,
  output LIOB33_X0Y83_IOB_X0Y84_OPAD,
  output LIOB33_X0Y85_IOB_X0Y85_OPAD,
  output LIOB33_X0Y85_IOB_X0Y86_OPAD,
  output LIOB33_X0Y87_IOB_X0Y87_OPAD,
  output LIOB33_X0Y87_IOB_X0Y88_OPAD,
  output LIOB33_X0Y89_IOB_X0Y89_OPAD,
  output LIOB33_X0Y89_IOB_X0Y90_OPAD,
  output LIOB33_X0Y91_IOB_X0Y91_OPAD,
  output LIOB33_X0Y91_IOB_X0Y92_OPAD,
  output LIOB33_X0Y93_IOB_X0Y93_OPAD,
  output LIOB33_X0Y93_IOB_X0Y94_OPAD,
  output LIOB33_X0Y95_IOB_X0Y95_OPAD,
  output LIOB33_X0Y95_IOB_X0Y96_OPAD,
  output LIOB33_X0Y97_IOB_X0Y97_OPAD,
  output LIOB33_X0Y97_IOB_X0Y98_OPAD,
  output RIOB33_SING_X105Y100_IOB_X1Y100_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_SING_X105Y50_IOB_X1Y50_OPAD,
  output RIOB33_SING_X105Y99_IOB_X1Y99_OPAD,
  output RIOB33_X105Y101_IOB_X1Y101_OPAD,
  output RIOB33_X105Y101_IOB_X1Y102_OPAD,
  output RIOB33_X105Y103_IOB_X1Y103_OPAD,
  output RIOB33_X105Y103_IOB_X1Y104_OPAD,
  output RIOB33_X105Y105_IOB_X1Y105_OPAD,
  output RIOB33_X105Y105_IOB_X1Y106_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD,
  output RIOB33_X105Y51_IOB_X1Y51_OPAD,
  output RIOB33_X105Y51_IOB_X1Y52_OPAD,
  output RIOB33_X105Y53_IOB_X1Y53_OPAD,
  output RIOB33_X105Y53_IOB_X1Y54_OPAD,
  output RIOB33_X105Y55_IOB_X1Y55_OPAD,
  output RIOB33_X105Y55_IOB_X1Y56_OPAD,
  output RIOB33_X105Y57_IOB_X1Y57_OPAD,
  output RIOB33_X105Y57_IOB_X1Y58_OPAD,
  output RIOB33_X105Y59_IOB_X1Y59_OPAD,
  output RIOB33_X105Y59_IOB_X1Y60_OPAD,
  output RIOB33_X105Y61_IOB_X1Y61_OPAD,
  output RIOB33_X105Y61_IOB_X1Y62_OPAD,
  output RIOB33_X105Y63_IOB_X1Y63_OPAD,
  output RIOB33_X105Y63_IOB_X1Y64_OPAD,
  output RIOB33_X105Y65_IOB_X1Y65_OPAD,
  output RIOB33_X105Y65_IOB_X1Y66_OPAD,
  output RIOB33_X105Y67_IOB_X1Y67_OPAD,
  output RIOB33_X105Y67_IOB_X1Y68_OPAD,
  output RIOB33_X105Y69_IOB_X1Y69_OPAD,
  output RIOB33_X105Y69_IOB_X1Y70_OPAD,
  output RIOB33_X105Y71_IOB_X1Y71_OPAD,
  output RIOB33_X105Y71_IOB_X1Y72_OPAD,
  output RIOB33_X105Y73_IOB_X1Y73_OPAD,
  output RIOB33_X105Y73_IOB_X1Y74_OPAD,
  output RIOB33_X105Y75_IOB_X1Y75_OPAD,
  output RIOB33_X105Y75_IOB_X1Y76_OPAD,
  output RIOB33_X105Y77_IOB_X1Y77_OPAD,
  output RIOB33_X105Y79_IOB_X1Y79_OPAD,
  output RIOB33_X105Y79_IOB_X1Y80_OPAD,
  output RIOB33_X105Y81_IOB_X1Y81_OPAD,
  output RIOB33_X105Y81_IOB_X1Y82_OPAD,
  output RIOB33_X105Y83_IOB_X1Y83_OPAD,
  output RIOB33_X105Y83_IOB_X1Y84_OPAD,
  output RIOB33_X105Y85_IOB_X1Y85_OPAD,
  output RIOB33_X105Y85_IOB_X1Y86_OPAD,
  output RIOB33_X105Y87_IOB_X1Y87_OPAD,
  output RIOB33_X105Y87_IOB_X1Y88_OPAD,
  output RIOB33_X105Y89_IOB_X1Y89_OPAD,
  output RIOB33_X105Y89_IOB_X1Y90_OPAD,
  output RIOB33_X105Y91_IOB_X1Y91_OPAD,
  output RIOB33_X105Y91_IOB_X1Y92_OPAD,
  output RIOB33_X105Y93_IOB_X1Y93_OPAD,
  output RIOB33_X105Y93_IOB_X1Y94_OPAD,
  output RIOB33_X105Y95_IOB_X1Y95_OPAD,
  output RIOB33_X105Y95_IOB_X1Y96_OPAD,
  output RIOB33_X105Y97_IOB_X1Y97_OPAD,
  output RIOB33_X105Y97_IOB_X1Y98_OPAD
  );
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A5Q;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_AMUX;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_AO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_AO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_AQ;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_A_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B5Q;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_BMUX;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_BO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_BO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_BQ;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_B_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_CLK;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_CO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_CO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_C_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_DO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_DO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_D_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X156Y111_SR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A5Q;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_AMUX;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_AO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_AO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_AQ;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_A_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B5Q;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_BMUX;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_BO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_BO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_BQ;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_B_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C5Q;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_CLK;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_CMUX;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_CO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_CO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_CQ;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_C_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D1;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D2;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D3;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D4;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_DMUX;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_DO5;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_DO6;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D_CY;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_D_XOR;
  wire [0:0] CLBLL_L_X100Y111_SLICE_X157Y111_SR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A5Q;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_AMUX;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_AO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_AO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_AQ;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_A_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_BO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_BO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_B_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_CLK;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_CO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_CO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_C_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_DO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_DO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_D_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X156Y112_SR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A5Q;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_AMUX;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_AO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_AO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_AQ;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_A_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_BO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_BO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_B_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_CLK;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_CO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_CO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_C_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D1;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D2;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D3;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D4;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_DO5;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_DO6;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D_CY;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_D_XOR;
  wire [0:0] CLBLL_L_X100Y112_SLICE_X157Y112_SR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A5Q;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_AMUX;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_AO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_AQ;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B5Q;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_BMUX;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_BO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_BQ;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C5Q;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CLK;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CMUX;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CQ;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_DO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_DO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_SR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A5Q;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_AMUX;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_AO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_AO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_AQ;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_BO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_BO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_CLK;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_CO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_CO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_DO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_DO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_SR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A5Q;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_AMUX;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_AO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_AO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_AQ;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_A_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B5Q;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_BMUX;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_BO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_BO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_BQ;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_B_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_CLK;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_CO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_CO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_C_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_DMUX;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_DO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_DO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_D_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X156Y114_SR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_AO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_AO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_A_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_BO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_BO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_B_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_CO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_CO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_C_XOR;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D1;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D2;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D3;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D4;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_DO5;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_DO6;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D_CY;
  wire [0:0] CLBLL_L_X100Y114_SLICE_X157Y114_D_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A5Q;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_AMUX;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_AO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_AO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_AQ;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_A_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B5Q;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_BMUX;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_BO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_BO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_BQ;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_B_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C5Q;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_CLK;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_CMUX;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_CO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_CO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_CQ;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_C_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_DO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_DO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_D_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X156Y115_SR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_AO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_AO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_AQ;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_A_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B5Q;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_BMUX;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_BO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_BO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_BQ;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_B_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_CLK;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_CO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_CO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_C_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D1;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D2;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D3;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D4;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_DMUX;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_DO5;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_DO6;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D_CY;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_D_XOR;
  wire [0:0] CLBLL_L_X100Y115_SLICE_X157Y115_SR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A5Q;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_AMUX;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_AO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_AO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_AQ;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_A_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B5Q;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_BMUX;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_BO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_BO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_BQ;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_B_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_CLK;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_CMUX;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_CO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_CO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_C_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_DO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_DO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_D_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X156Y116_SR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A5Q;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_AMUX;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_AO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_AO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_AQ;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_A_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B5Q;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_BMUX;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_BO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_BO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_BQ;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_B_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_CLK;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_CO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_CO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_C_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D1;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D2;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D3;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D4;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_DO5;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_DO6;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D_CY;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_D_XOR;
  wire [0:0] CLBLL_L_X100Y116_SLICE_X157Y116_SR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A5Q;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_AMUX;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_AO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_AO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_AQ;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_A_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B5Q;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_BMUX;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_BO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_BO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_BQ;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_B_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_CLK;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_CMUX;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_CO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_CO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_C_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_DO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_DO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_D_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X156Y117_SR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A5Q;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_AMUX;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_AO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_AO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_AQ;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_A_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B5Q;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_BMUX;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_BO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_BO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_BQ;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_B_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_CLK;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_CO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_CO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_C_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D1;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D2;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D3;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D4;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_DO5;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_DO6;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D_CY;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_D_XOR;
  wire [0:0] CLBLL_L_X100Y117_SLICE_X157Y117_SR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A5Q;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_AMUX;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_AO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_AO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_AQ;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_A_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B5Q;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_BMUX;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_BO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_BO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_BQ;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_B_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_CLK;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_CO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_CO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_C_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_DO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_DO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_D_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X156Y118_SR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A5Q;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_AMUX;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_AO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_AO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_AQ;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_A_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B5Q;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_BMUX;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_BO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_BO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_BQ;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_B_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C5Q;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_CLK;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_CMUX;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_CO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_CO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_CQ;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_C_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D1;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D2;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D3;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D4;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_DO5;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_DO6;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D_CY;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_D_XOR;
  wire [0:0] CLBLL_L_X100Y118_SLICE_X157Y118_SR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_AO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_AO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_AQ;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_A_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B5Q;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_BMUX;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_BO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_BO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_BQ;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_B_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_CLK;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_CO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_CO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_C_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_DO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_DO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_D_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X156Y119_SR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A5Q;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_AMUX;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_AO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_AO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_AQ;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_AX;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_A_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_BMUX;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_BO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_BO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_B_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C5Q;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_CLK;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_CMUX;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_CO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_CO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_CQ;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_C_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D1;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D2;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D3;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D4;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_DO5;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_DO6;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D_CY;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_D_XOR;
  wire [0:0] CLBLL_L_X100Y119_SLICE_X157Y119_SR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_AO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_AO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_AQ;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_A_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_BO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_BO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_B_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_CLK;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_CO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_CO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_C_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_DO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_DO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_D_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X156Y120_SR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A5Q;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_AMUX;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_AO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_AO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_AQ;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_A_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_BO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_BO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_BQ;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_B_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_CLK;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_CO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_CO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_C_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D1;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D2;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D3;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D4;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_DO5;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_DO6;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D_CY;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_D_XOR;
  wire [0:0] CLBLL_L_X100Y120_SLICE_X157Y120_SR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A5Q;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_AMUX;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_AO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_AQ;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_BO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_BQ;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C5Q;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CLK;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CMUX;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CQ;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_DO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_DO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_SR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_AO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_AO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_AQ;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_BO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_BO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_BQ;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C5Q;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CLK;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CMUX;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CQ;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_DO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_DO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_SR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A5Q;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_AMUX;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_AO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_AO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_AQ;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_A_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_BO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_BO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_B_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_CLK;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_CO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_CO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_C_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_DO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_DO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_D_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X156Y122_SR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A5Q;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_AMUX;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_AO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_AO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_AQ;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_A_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B5Q;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_BMUX;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_BO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_BO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_BQ;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_B_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C5Q;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_CLK;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_CMUX;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_CO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_CO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_CQ;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_C_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D1;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D2;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D3;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D4;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_DO5;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_DO6;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D_CY;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_D_XOR;
  wire [0:0] CLBLL_L_X100Y122_SLICE_X157Y122_SR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A5Q;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AMUX;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AQ;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B5Q;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BMUX;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BQ;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_CLK;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_CO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_CO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_DO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_DO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_SR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A5Q;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_AMUX;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_AO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_AO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_AQ;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_BO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_BO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_CLK;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_CO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_CO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_DO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_DO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_SR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_AMUX;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_AO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_AO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_AQ;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_A_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B5Q;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_BMUX;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_BO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_BO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_BQ;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_B_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_CLK;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_CO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_CO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_C_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_DO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_DO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_D_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X156Y124_SR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A5Q;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_AMUX;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_AO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_AO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_AQ;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_A_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B5Q;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_BMUX;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_BO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_BO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_BQ;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_B_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_CLK;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_CO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_CO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_C_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D1;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D2;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D3;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D4;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_DO5;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_DO6;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D_CY;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_D_XOR;
  wire [0:0] CLBLL_L_X100Y124_SLICE_X157Y124_SR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_AO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_AO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_AQ;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_A_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B5Q;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_BMUX;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_BO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_BO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_BQ;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_B_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_CLK;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_CO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_CO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_C_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_DO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_DO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_D_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X156Y125_SR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A5Q;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_AMUX;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_AO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_AO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_AQ;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_A_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B5Q;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_BMUX;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_BO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_BO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_BQ;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_B_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C5Q;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_CLK;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_CMUX;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_CO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_CO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_CQ;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_C_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D1;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D2;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D3;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D4;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_DO5;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_DO6;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_DQ;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D_CY;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_D_XOR;
  wire [0:0] CLBLL_L_X100Y125_SLICE_X157Y125_SR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A5Q;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_AMUX;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_AO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_AO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_AQ;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_A_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B5Q;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_BMUX;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_BO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_BO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_BQ;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_B_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_CLK;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_CMUX;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_CO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_CO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_C_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_DO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_DO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_D_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X156Y126_SR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A5Q;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_AMUX;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_AO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_AO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_AQ;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_A_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_BO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_BO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_BQ;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_B_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_CLK;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_CO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_CO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_CQ;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_C_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D1;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D2;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D3;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D4;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_DO5;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_DO6;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D_CY;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_D_XOR;
  wire [0:0] CLBLL_L_X100Y126_SLICE_X157Y126_SR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A5Q;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_AMUX;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_AO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_AO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_AQ;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_A_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B5Q;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_BMUX;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_BO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_BO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_BQ;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_B_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_CLK;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_CO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_CO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_C_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_DO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_DO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_D_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X156Y127_SR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_AO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_AO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_AQ;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_A_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B5Q;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_BMUX;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_BO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_BO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_BQ;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_B_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_CLK;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_CO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_CO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_C_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D1;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D2;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D3;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D4;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_DO5;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_DO6;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D_CY;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_D_XOR;
  wire [0:0] CLBLL_L_X100Y127_SLICE_X157Y127_SR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A5Q;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_AMUX;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_AO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_AO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_AQ;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_A_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_BO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_BO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_BQ;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_B_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_CLK;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_CO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_CO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_C_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_DO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_DO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_D_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X156Y128_SR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_AO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_AO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_A_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_BO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_BO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_B_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_CO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_CO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_C_XOR;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D1;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D2;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D3;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D4;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_DO5;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_DO6;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D_CY;
  wire [0:0] CLBLL_L_X100Y128_SLICE_X157Y128_D_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_AO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_AO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_AQ;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_A_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_BO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_BO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_B_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_CLK;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_CO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_CO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_C_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_DO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_DO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_D_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X156Y129_SR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A5Q;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_AMUX;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_AO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_AO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_AQ;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_A_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_BO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_BO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_B_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_CLK;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_CO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_CO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_C_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D1;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D2;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D3;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D4;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_DO5;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_DO6;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D_CY;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_D_XOR;
  wire [0:0] CLBLL_L_X100Y129_SLICE_X157Y129_SR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_AO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_AO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_AQ;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_A_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_BO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_BO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_B_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_CLK;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_CO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_CO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_C_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_DO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_DO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_D_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X156Y130_SR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_AO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_AO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_A_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_BO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_BO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_B_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_CO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_CO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_C_XOR;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D1;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D2;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D3;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D4;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_DO5;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_DO6;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D_CY;
  wire [0:0] CLBLL_L_X100Y130_SLICE_X157Y130_D_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A5Q;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_AMUX;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_AO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_AO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_AQ;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_A_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_BO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_BO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_B_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_CLK;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_CO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_CO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_C_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_DO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_DO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_D_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X156Y133_SR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_AO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_AO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_A_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_BO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_BO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_B_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_CO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_CO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_C_XOR;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D1;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D2;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D3;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D4;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_DO5;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_DO6;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D_CY;
  wire [0:0] CLBLL_L_X100Y133_SLICE_X157Y133_D_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A5Q;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_AMUX;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_AO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_AO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_AQ;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_A_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B5Q;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_BMUX;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_BO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_BO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_BQ;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_B_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_CLK;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_CO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_CO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_C_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_DO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_DO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_D_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X156Y134_SR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_AO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_AO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_A_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_BO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_BO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_B_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_CO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_CO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_C_XOR;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D1;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D2;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D3;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D4;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_DO5;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_DO6;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D_CY;
  wire [0:0] CLBLL_L_X100Y134_SLICE_X157Y134_D_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CLK;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_SR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B5Q;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CLK;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_DO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_DO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_SR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CLK;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_SR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CLK;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_DO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_DO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_SR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A5Q;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_AMUX;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_AO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_AO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_AQ;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_BO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_BO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_CLK;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_CO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_CO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_DO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_DO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_SR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A5Q;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AMUX;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B5Q;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_BMUX;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_BO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_BO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_BQ;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CLK;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CMUX;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_DO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_DO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_SR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_AMUX;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_AO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B5Q;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_BMUX;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_BO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_BO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_BQ;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C5Q;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CLK;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CMUX;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CQ;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_DO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_DO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_SR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A5Q;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AMUX;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_BO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_BO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_CLK;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_CO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_CO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_DO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_DO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_SR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A5Q;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B5Q;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_BMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_BO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_BO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_BQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CLK;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_DO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_DO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_SR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B5Q;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C5Q;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CLK;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_DO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_SR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_AMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_AO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_AO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_AQ;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_AX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_A_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B5Q;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_BMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_BO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_BO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_BQ;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_B_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C5Q;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_CLK;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_CMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_CO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_CO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_CQ;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_C_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_DO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_DO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_D_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X160Y116_SR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A5Q;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_AMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_AO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_AO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_AQ;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_A_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B5Q;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_BMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_BO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_BO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_BQ;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_B_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_CLK;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_CMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_CO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_CO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_CQ;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_CX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_C_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D1;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D2;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D3;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D4;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_DMUX;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_DO5;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_DO6;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D_CY;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_D_XOR;
  wire [0:0] CLBLL_L_X102Y116_SLICE_X161Y116_SR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_AO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_AO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_AQ;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_A_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B5Q;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_BMUX;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_BO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_BO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_BQ;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_B_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_CLK;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_CO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_CO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_C_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_DO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_DO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_D_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X160Y117_SR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A5Q;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_AMUX;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_AO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_AO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_AQ;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_A_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B5Q;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_BMUX;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_BO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_BO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_BQ;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_B_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C5Q;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_CLK;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_CMUX;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_CO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_CO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_CQ;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_C_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D1;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D2;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D3;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D4;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D5Q;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_DMUX;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_DO5;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_DO6;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_DQ;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D_CY;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_D_XOR;
  wire [0:0] CLBLL_L_X102Y117_SLICE_X161Y117_SR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_AMUX;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_AO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_AO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_A_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_BO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_BO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_B_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_CO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_CO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_C_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_DO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_DO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X160Y118_D_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_AO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_AO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_A_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_BO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_BO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_B_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_CO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_CO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_C_XOR;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D1;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D2;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D3;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D4;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_DO5;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_DO6;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D_CY;
  wire [0:0] CLBLL_L_X102Y118_SLICE_X161Y118_D_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A5Q;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_AMUX;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_AO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_AO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_AQ;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_A_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B5Q;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_BMUX;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_BO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_BO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_BQ;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_B_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_CLK;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_CO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_CO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_C_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_DO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_DO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_D_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X160Y119_SR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_AO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_AO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_AQ;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_A_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B5Q;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_BMUX;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_BO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_BO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_BQ;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_B_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_CLK;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_CO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_CO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_C_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D1;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D2;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D3;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D4;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_DO5;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_DO6;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D_CY;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_D_XOR;
  wire [0:0] CLBLL_L_X102Y119_SLICE_X161Y119_SR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_AO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_AO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_AQ;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_A_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B5Q;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_BMUX;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_BO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_BO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_BQ;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_B_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C5Q;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_CLK;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_CMUX;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_CO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_CO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_CQ;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_C_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D5Q;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_DMUX;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_DO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_DO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_DQ;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_D_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X160Y120_SR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_AO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_AO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_AQ;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_A_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B5Q;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_BMUX;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_BO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_BO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_BQ;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_B_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_CLK;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_CO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_CO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_C_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D1;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D2;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D3;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D4;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_DMUX;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_DO5;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_DO6;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D_CY;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_D_XOR;
  wire [0:0] CLBLL_L_X102Y120_SLICE_X161Y120_SR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_AO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_AO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_AQ;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_A_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_BO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_BO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_B_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_CLK;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_CO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_CO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_C_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_DO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_DO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_D_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X160Y121_SR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A5Q;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_AMUX;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_AO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_AO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_AQ;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_A_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B5Q;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_BMUX;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_BO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_BO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_BQ;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_B_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C5Q;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_CLK;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_CMUX;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_CO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_CO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_CQ;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_C_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D1;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D2;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D3;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D4;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_DO5;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_DO6;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D_CY;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_D_XOR;
  wire [0:0] CLBLL_L_X102Y121_SLICE_X161Y121_SR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A5Q;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_AMUX;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_AO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_AO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_AQ;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_A_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B5Q;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_BMUX;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_BO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_BO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_BQ;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_B_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C5Q;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_CLK;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_CMUX;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_CO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_CO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_CQ;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_C_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_DO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_DO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_D_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X160Y122_SR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A5Q;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_AMUX;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_AO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_AO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_AQ;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_A_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B5Q;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_BMUX;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_BO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_BO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_BQ;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_B_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C5Q;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_CLK;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_CMUX;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_CO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_CO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_CQ;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_C_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D1;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D2;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D3;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D4;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_DO5;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_DO6;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D_CY;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_D_XOR;
  wire [0:0] CLBLL_L_X102Y122_SLICE_X161Y122_SR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_AO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_AO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_AQ;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_A_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B5Q;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_BMUX;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_BO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_BO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_BQ;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_B_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_CLK;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_CO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_CO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_C_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_DO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_DO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_D_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X160Y123_SR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A5Q;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_AMUX;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_AO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_AO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_AQ;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_A_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_BO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_BO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_B_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_CLK;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_CO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_CO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_C_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D1;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D2;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D3;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D4;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_DMUX;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_DO5;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_DO6;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D_CY;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_D_XOR;
  wire [0:0] CLBLL_L_X102Y123_SLICE_X161Y123_SR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A5Q;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_AMUX;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_AO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_AO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_AQ;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_A_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_BO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_BO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_BQ;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_B_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C5Q;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_CLK;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_CMUX;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_CO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_CO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_CQ;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_C_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D5Q;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_DMUX;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_DO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_DO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_DQ;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_D_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X160Y124_SR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A5Q;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_AMUX;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_AO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_AO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_AQ;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_A_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B5Q;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_BMUX;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_BO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_BO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_BQ;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_B_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_CLK;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_CO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_CO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_C_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D1;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D2;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D3;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D4;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_DO5;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_DO6;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D_CY;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_D_XOR;
  wire [0:0] CLBLL_L_X102Y124_SLICE_X161Y124_SR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_AO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_AO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_AQ;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_A_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B5Q;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_BMUX;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_BO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_BO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_BQ;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_B_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_CLK;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_CO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_CO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_C_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_DO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_DO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_D_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X160Y125_SR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_AO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_AQ;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_A_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B5Q;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_BMUX;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_BO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_BQ;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_B_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C5Q;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CLK;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CMUX;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_CQ;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_C_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D1;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D2;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D3;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D4;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_DMUX;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_DO5;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D_CY;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_D_XOR;
  wire [0:0] CLBLL_L_X102Y125_SLICE_X161Y125_SR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A5Q;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_AMUX;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_AO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_AO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_AQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_A_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_BO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_BO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_BQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_B_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C5Q;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_CLK;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_CMUX;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_CO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_CO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_CQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_C_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_DO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_DO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_D_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X160Y126_SR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A5Q;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_AMUX;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_AO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_AO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_AQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_A_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B5Q;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_BMUX;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_BO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_BO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_BQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_B_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C5Q;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_CLK;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_CMUX;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_CO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_CO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_CQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_C_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D1;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D2;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D3;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D4;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D5Q;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_DMUX;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_DO5;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_DO6;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_DQ;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D_CY;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_D_XOR;
  wire [0:0] CLBLL_L_X102Y126_SLICE_X161Y126_SR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A5Q;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_AMUX;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_AO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_AO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_AQ;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_A_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_BO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_BO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_BQ;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_B_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C5Q;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_CLK;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_CMUX;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_CO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_CO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_CQ;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_C_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_DO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_DO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_D_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X160Y127_SR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A5Q;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_AMUX;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_AO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_AO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_AQ;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_A_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B5Q;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_BMUX;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_BO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_BO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_BQ;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_B_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_CLK;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_CO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_CO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_C_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D1;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D2;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D3;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D4;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_DO5;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_DO6;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D_CY;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_D_XOR;
  wire [0:0] CLBLL_L_X102Y127_SLICE_X161Y127_SR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_AO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_AO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_A_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_BO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_BO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_B_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_CO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_CO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_C_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_DO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_DO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X160Y128_D_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_AO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_AO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_AQ;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_A_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B5Q;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_BMUX;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_BO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_BO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_BQ;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_B_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_CLK;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_CO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_CO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_C_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D1;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D2;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D3;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D4;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_DO5;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_DO6;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D_CY;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_D_XOR;
  wire [0:0] CLBLL_L_X102Y128_SLICE_X161Y128_SR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A5Q;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_AMUX;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_AO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_AO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_AQ;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_A_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_BO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_BO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_BQ;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_B_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C5Q;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_CLK;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_CMUX;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_CO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_CO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_CQ;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_C_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_DO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_DO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_D_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X160Y129_SR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_AO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_AO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_AQ;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_A_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_BO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_BO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_B_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_CLK;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_CO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_CO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_C_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D1;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D2;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D3;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D4;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_DO5;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_DO6;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D_CY;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_D_XOR;
  wire [0:0] CLBLL_L_X102Y129_SLICE_X161Y129_SR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A5Q;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_AMUX;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_AO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_AO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_AQ;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_A_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B5Q;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_BMUX;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_BO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_BO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_BQ;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_B_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_CLK;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_CMUX;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_CO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_CO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_C_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_DO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_DO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_D_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X160Y130_SR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A5Q;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_AMUX;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_AO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_AO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_AQ;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_A_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_BO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_BO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_BQ;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_B_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_CLK;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_CO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_CO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_C_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D1;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D2;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D3;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D4;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_DO5;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_DO6;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D_CY;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_D_XOR;
  wire [0:0] CLBLL_L_X102Y130_SLICE_X161Y130_SR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_AO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_AO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_AQ;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_A_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B5Q;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_BMUX;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_BO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_BO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_BQ;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_B_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_CLK;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_CO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_CO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_C_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_DO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_DO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_D_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X160Y131_SR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_AO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_AO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_A_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_BO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_BO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_B_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_CO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_CO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_C_XOR;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D1;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D2;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D3;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D4;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_DO5;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_DO6;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D_CY;
  wire [0:0] CLBLL_L_X102Y131_SLICE_X161Y131_D_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A5Q;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_AMUX;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_AO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_AO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_AQ;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_A_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_BO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_BO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_B_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_CLK;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_CO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_CO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_C_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_DO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_DO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_D_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X160Y134_SR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_AO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_AO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_A_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_BO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_BO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_B_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_CO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_CO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_C_XOR;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D1;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D2;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D3;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D4;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_DO5;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_DO6;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D_CY;
  wire [0:0] CLBLL_L_X102Y134_SLICE_X161Y134_D_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_AO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_AO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_AQ;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_A_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_BO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_BO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_B_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_CLK;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_CO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_CO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_C_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_DO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_DO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_D_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X160Y135_SR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_AO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_AO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_A_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_BO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_BO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_B_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_CO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_CO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_C_XOR;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D1;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D2;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D3;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D4;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_DO5;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_DO6;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D_CY;
  wire [0:0] CLBLL_L_X102Y135_SLICE_X161Y135_D_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_AO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_AO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_AQ;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_A_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B5Q;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_BMUX;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_BO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_BO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_BQ;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_B_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_CLK;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_CO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_CO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_C_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_DO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_DO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_D_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X160Y136_SR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_AO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_AO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_A_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_BO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_BO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_B_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_CO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_CO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_C_XOR;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D1;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D2;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D3;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D4;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_DO5;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_DO6;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D_CY;
  wire [0:0] CLBLL_L_X102Y136_SLICE_X161Y136_D_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_AO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_AO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_AQ;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_A_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B5Q;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_BMUX;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_BO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_BO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_BQ;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_B_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_CLK;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_CO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_CO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_C_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_DO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_DO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_D_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X138Y118_SR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_AO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_AO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_AQ;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_A_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_BO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_BO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_B_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_CLK;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_CO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_CO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_C_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D1;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D2;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D3;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D4;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_DO5;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_DO6;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D_CY;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_D_XOR;
  wire [0:0] CLBLL_R_X87Y118_SLICE_X139Y118_SR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A5Q;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_AMUX;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_AO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_AO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_AQ;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_A_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_BO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_BO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_B_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_CLK;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_CO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_CO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_C_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_DO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_DO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_D_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X142Y113_SR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A5Q;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_AMUX;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_AO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_AO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_AQ;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_A_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B5Q;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_BMUX;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_BO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_BO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_BQ;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_B_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C5Q;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_CLK;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_CMUX;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_CO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_CO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_CQ;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_C_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D1;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D2;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D3;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D4;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_DO5;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_DO6;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D_CY;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_D_XOR;
  wire [0:0] CLBLM_L_X90Y113_SLICE_X143Y113_SR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A5Q;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_AMUX;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_AO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_AO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_AQ;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_A_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B5Q;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_BMUX;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_BO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_BO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_BQ;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_B_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C5Q;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_CLK;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_CMUX;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_CO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_CO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_CQ;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_C_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_DO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_DO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_D_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X142Y114_SR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A5Q;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_AMUX;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_AO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_AO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_AQ;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_A_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B5Q;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_BMUX;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_BO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_BO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_BQ;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_B_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_CLK;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_CMUX;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_CO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_CO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_C_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D1;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D2;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D3;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D4;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_DO5;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_DO6;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D_CY;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_D_XOR;
  wire [0:0] CLBLM_L_X90Y114_SLICE_X143Y114_SR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A5Q;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_AMUX;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_AO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_AO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_AQ;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_A_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_BO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_BO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_BQ;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_B_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_CLK;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_CO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_CO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_C_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_DO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_DO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_D_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X142Y115_SR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A5Q;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_AMUX;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_AO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_AO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_AQ;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_A_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B5Q;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_BMUX;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_BO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_BO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_BQ;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_B_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C5Q;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_CLK;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_CMUX;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_CO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_CO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_CQ;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_C_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D1;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D2;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D3;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D4;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_DMUX;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_DO5;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_DO6;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D_CY;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_D_XOR;
  wire [0:0] CLBLM_L_X90Y115_SLICE_X143Y115_SR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A5Q;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_AMUX;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_AO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_AO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_AQ;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_A_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_BO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_BO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_BQ;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_B_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C5Q;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_CLK;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_CMUX;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_CO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_CO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_CQ;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_C_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_DO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_DO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_D_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X142Y116_SR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A5Q;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_AMUX;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_AO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_AO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_AQ;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_A_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B5Q;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_BMUX;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_BO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_BO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_BQ;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_B_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C5Q;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_CLK;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_CMUX;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_CO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_CO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_CQ;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_C_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D1;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D2;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D3;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D4;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_DO5;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_DO6;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D_CY;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_D_XOR;
  wire [0:0] CLBLM_L_X90Y116_SLICE_X143Y116_SR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A5Q;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_AMUX;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_AO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_AO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_AQ;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_AX;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_A_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_BMUX;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_BO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_BO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_B_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C5Q;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_CLK;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_CMUX;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_CO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_CO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_CQ;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_C_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_DO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_DO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_D_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X142Y117_SR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A5Q;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_AMUX;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_AO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_AO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_AQ;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_A_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B5Q;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_BMUX;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_BO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_BO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_BQ;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_B_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_CLK;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_CO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_CO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_C_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D1;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D2;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D3;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D4;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_DO5;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_DO6;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D_CY;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_D_XOR;
  wire [0:0] CLBLM_L_X90Y117_SLICE_X143Y117_SR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A5Q;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_AMUX;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_AO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_AO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_AQ;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_A_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B5Q;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_BMUX;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_BO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_BO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_BQ;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_B_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_CLK;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_CO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_CO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_C_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_DMUX;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_DO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_DO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_D_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X142Y118_SR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A5Q;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_AMUX;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_AO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_AO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_AQ;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_A_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B5Q;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_BMUX;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_BO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_BO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_BQ;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_B_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_CLK;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_CO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_CO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_C_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D1;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D2;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D3;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D4;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_DMUX;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_DO5;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_DO6;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D_CY;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_D_XOR;
  wire [0:0] CLBLM_L_X90Y118_SLICE_X143Y118_SR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_AMUX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_AO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_AO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_A_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B5Q;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_BMUX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_BO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_BO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_BQ;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_B_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C5Q;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_CLK;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_CMUX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_CO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_CO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_CQ;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_C_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_DO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_DO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_D_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X142Y119_SR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_AMUX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_AO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_AO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_AQ;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_AX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_A_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B5Q;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_BMUX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_BO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_BO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_BQ;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_B_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_CLK;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_CO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_CO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_CQ;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_CX;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_C_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D1;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D2;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D3;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D4;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_DO5;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_DO6;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D_CY;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_D_XOR;
  wire [0:0] CLBLM_L_X90Y119_SLICE_X143Y119_SR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A5Q;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_AMUX;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_AO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_AO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_AQ;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_A_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B5Q;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_BMUX;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_BO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_BO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_BQ;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_BX;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_B_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_CLK;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_CMUX;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_CO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_CO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_C_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_DO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_DO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_D_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X142Y120_SR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A5Q;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_AMUX;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_AO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_AO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_AQ;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_A_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_BO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_BO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_BQ;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_B_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C5Q;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_CLK;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_CMUX;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_CO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_CO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_CQ;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_C_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D1;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D2;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D3;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D4;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_DO5;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_DO6;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D_CY;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_D_XOR;
  wire [0:0] CLBLM_L_X90Y120_SLICE_X143Y120_SR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A5Q;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_AMUX;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_AO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_AO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_AQ;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_A_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_BO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_BO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_B_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_CLK;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_CO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_CO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_C_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_DO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_DO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_D_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X142Y121_SR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A5Q;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_AMUX;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_AO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_AO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_AQ;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_AX;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_A_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_BMUX;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_BO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_BO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_B_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C5Q;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_CLK;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_CMUX;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_CO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_CO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_CQ;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_C_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D1;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D2;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D3;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D4;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_DO5;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_DO6;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D_CY;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_D_XOR;
  wire [0:0] CLBLM_L_X90Y121_SLICE_X143Y121_SR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A5Q;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_AMUX;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_AO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_AO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_AQ;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_A_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_BO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_BO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_BQ;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_B_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_CLK;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_CO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_CO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_C_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_DO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_DO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_D_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X142Y122_SR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A5Q;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_AMUX;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_AO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_AO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_AQ;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_AX;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_A_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_BMUX;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_BO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_BO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_B_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C5Q;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_CLK;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_CMUX;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_CO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_CO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_CQ;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_C_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D1;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D2;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D3;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D4;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_DO5;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_DO6;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D_CY;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_D_XOR;
  wire [0:0] CLBLM_L_X90Y122_SLICE_X143Y122_SR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A5Q;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_AMUX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_AO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_AO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_AQ;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_A_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B5Q;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_BMUX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_BO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_BO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_BQ;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_B_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C5Q;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_CLK;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_CMUX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_CO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_CO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_CQ;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_C_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_DO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_DO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_D_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X142Y123_SR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A5Q;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_AMUX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_AO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_AO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_AQ;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_AX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_A_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_BMUX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_BO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_BO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_B_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C5Q;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_CLK;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_CMUX;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_CO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_CO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_CQ;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_C_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D1;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D2;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D3;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D4;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_DO5;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_DO6;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D_CY;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_D_XOR;
  wire [0:0] CLBLM_L_X90Y123_SLICE_X143Y123_SR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A5Q;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_AMUX;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_AO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_AO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_AQ;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_AX;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_A_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_BMUX;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_BO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_BO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_B_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C5Q;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_CLK;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_CMUX;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_CO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_CO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_CQ;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_C_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_DO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_DO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_D_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X142Y124_SR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_AO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_AO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_AQ;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_A_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B5Q;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_BMUX;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_BO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_BO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_BQ;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_B_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C5Q;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_CLK;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_CMUX;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_CO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_CO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_CQ;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_C_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D1;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D2;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D3;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D4;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_DO5;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_DO6;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D_CY;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_D_XOR;
  wire [0:0] CLBLM_L_X90Y124_SLICE_X143Y124_SR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A5Q;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_AMUX;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_AO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_AO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_AQ;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_A_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_BO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_BO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_B_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_CLK;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_CO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_CO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_C_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_DO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_DO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_D_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X142Y125_SR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A5Q;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_AMUX;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_AO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_AO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_AQ;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_A_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B5Q;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_BMUX;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_BO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_BO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_BQ;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_B_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_CLK;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_CO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_CO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_CQ;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_C_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D1;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D2;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D3;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D4;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_DO5;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_DO6;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_DQ;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D_CY;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_D_XOR;
  wire [0:0] CLBLM_L_X90Y125_SLICE_X143Y125_SR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_AO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_AO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_AQ;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_A_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B5Q;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_BMUX;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_BO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_BO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_BQ;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_B_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C5Q;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_CLK;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_CMUX;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_CO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_CO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_CQ;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_C_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_DO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_DO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_D_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X142Y126_SR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A5Q;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_AMUX;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_AO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_AO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_AQ;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_AX;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_A_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_BMUX;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_BO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_BO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_B_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C5Q;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_CLK;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_CMUX;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_CO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_CO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_CQ;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_C_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D1;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D2;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D3;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D4;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_DO5;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_DO6;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D_CY;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_D_XOR;
  wire [0:0] CLBLM_L_X90Y126_SLICE_X143Y126_SR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_AMUX;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_AO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_AO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_AQ;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_A_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B5Q;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_BMUX;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_BO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_BO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_BQ;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_B_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_CLK;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_CO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_CO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_C_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_DO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_DO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_D_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X142Y128_SR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A5Q;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_AMUX;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_AO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_AO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_AQ;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_A_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_BO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_BO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_BQ;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_B_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_CLK;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_CO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_CO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_CQ;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_C_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D1;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D2;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D3;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D4;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D5Q;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_DMUX;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_DO5;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_DO6;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_DQ;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D_CY;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_D_XOR;
  wire [0:0] CLBLM_L_X90Y128_SLICE_X143Y128_SR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A5Q;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_AMUX;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_AO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_AO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_AQ;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_AX;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_A_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_BMUX;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_BO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_BO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_B_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C5Q;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_CLK;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_CMUX;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_CO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_CO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_CQ;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_C_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_DO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_DO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_D_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X142Y129_SR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_AO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_AO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_A_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_BO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_BO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_B_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_CO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_CO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_C_XOR;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D1;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D2;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D3;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D4;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_DO5;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_DO6;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D_CY;
  wire [0:0] CLBLM_L_X90Y129_SLICE_X143Y129_D_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A5Q;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_AMUX;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_AO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_AO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_AQ;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_A_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B5Q;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_BMUX;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_BO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_BO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_BQ;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_BX;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_B_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_CLK;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_CMUX;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_CO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_CO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_C_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_DO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_DO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_D_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X142Y130_SR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_AO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_AO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_A_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_BO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_BO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_B_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_CO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_CO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_C_XOR;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D1;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D2;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D3;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D4;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_DO5;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_DO6;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D_CY;
  wire [0:0] CLBLM_L_X90Y130_SLICE_X143Y130_D_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A5Q;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_AMUX;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_AO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_AO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_AQ;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_AX;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_A_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_BMUX;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_BO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_BO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_B_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C5Q;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_CLK;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_CMUX;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_CO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_CO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_CQ;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_C_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_DO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_DO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_D_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X142Y131_SR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_AO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_AO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_A_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_BO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_BO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_B_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_CO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_CO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_C_XOR;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D1;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D2;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D3;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D4;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_DO5;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_DO6;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D_CY;
  wire [0:0] CLBLM_L_X90Y131_SLICE_X143Y131_D_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_AO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_AO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_A_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_BO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_BO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_B_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_CO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_CO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_C_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_DO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_DO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X144Y112_D_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A5Q;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_AMUX;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_AO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_AO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_AQ;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_A_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B5Q;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_BMUX;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_BO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_BO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_BQ;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_B_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_CLK;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_CO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_CO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_C_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D1;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D2;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D3;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D4;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_DO5;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_DO6;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D_CY;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_D_XOR;
  wire [0:0] CLBLM_L_X92Y112_SLICE_X145Y112_SR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A5Q;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_AMUX;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_AO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_AO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_AQ;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_A_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B5Q;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_BMUX;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_BO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_BO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_BQ;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_B_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_CLK;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_CO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_CO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_C_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_DO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_DO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_D_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X144Y113_SR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A5Q;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_AMUX;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_AO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_AO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_AQ;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_A_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B5Q;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_BMUX;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_BO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_BO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_BQ;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_B_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_CLK;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_CO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_CO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_C_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D1;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D2;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D3;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D4;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_DO5;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_DO6;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D_CY;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_D_XOR;
  wire [0:0] CLBLM_L_X92Y113_SLICE_X145Y113_SR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A5Q;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_AMUX;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_AO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_AO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_AQ;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_A_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B5Q;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_BMUX;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_BO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_BO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_BQ;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_B_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_CLK;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_CO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_CO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_C_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_DO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_DO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_D_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X144Y114_SR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A5Q;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_AMUX;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_AO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_AO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_AQ;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_A_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_BO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_BO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_B_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_CLK;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_CO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_CO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_C_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D1;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D2;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D3;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D4;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_DO5;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_DO6;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D_CY;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_D_XOR;
  wire [0:0] CLBLM_L_X92Y114_SLICE_X145Y114_SR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_AO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_AO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_A_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_BO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_BO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_B_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_CO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_CO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_C_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_DO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_DO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X144Y115_D_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A5Q;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_AMUX;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_AO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_AO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_AQ;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_A_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B5Q;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_BMUX;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_BO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_BO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_BQ;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_B_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_CLK;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_CO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_CO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_C_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D1;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D2;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D3;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D4;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_DO5;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_DO6;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D_CY;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_D_XOR;
  wire [0:0] CLBLM_L_X92Y115_SLICE_X145Y115_SR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A5Q;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_AMUX;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_AO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_AO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_AQ;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_A_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B5Q;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_BMUX;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_BO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_BO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_BQ;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_B_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_CLK;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_CO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_CO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_C_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_DO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_DO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_D_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X144Y116_SR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A5Q;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_AMUX;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_AO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_AO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_AQ;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_A_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B5Q;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_BMUX;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_BO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_BO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_BQ;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_B_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_CLK;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_CO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_CO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_C_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D1;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D2;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D3;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D4;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_DO5;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_DO6;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D_CY;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_D_XOR;
  wire [0:0] CLBLM_L_X92Y116_SLICE_X145Y116_SR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A5Q;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_AMUX;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_AO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_AO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_AQ;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_A_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_BO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_BO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_B_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_CLK;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_CO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_CO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_C_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_DO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_DO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_D_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X144Y118_SR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_AO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_AO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_A_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_BO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_BO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_B_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_CO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_CO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_C_XOR;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D1;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D2;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D3;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D4;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_DO5;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_DO6;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D_CY;
  wire [0:0] CLBLM_L_X92Y118_SLICE_X145Y118_D_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A5Q;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_AMUX;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_AO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_AO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_AQ;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_AX;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_A_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_BMUX;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_BO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_BO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_B_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C5Q;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_CLK;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_CMUX;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_CO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_CO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_CQ;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_C_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_DO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_DO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_D_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X144Y119_SR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A5Q;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_AMUX;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_AO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_AO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_AQ;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_A_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B5Q;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_BMUX;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_BO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_BO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_BQ;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_B_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_CLK;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_CO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_CO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_C_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D1;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D2;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D3;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D4;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_DO5;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_DO6;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D_CY;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_D_XOR;
  wire [0:0] CLBLM_L_X92Y119_SLICE_X145Y119_SR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A5Q;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_AMUX;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_AO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_AO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_AQ;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_A_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B5Q;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_BMUX;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_BO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_BO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_BQ;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_B_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_CLK;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_CO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_CO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_C_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_DO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_DO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_D_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X144Y120_SR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A5Q;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_AMUX;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_AO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_AO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_AQ;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_AX;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_A_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_BMUX;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_BO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_BO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_B_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C5Q;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_CLK;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_CMUX;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_CO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_CO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_CQ;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_C_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D1;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D2;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D3;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D4;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_DO5;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_DO6;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D_CY;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_D_XOR;
  wire [0:0] CLBLM_L_X92Y120_SLICE_X145Y120_SR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A5Q;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_AMUX;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_AO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_AO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_AQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_A_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_BO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_BO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_BQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_B_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_CLK;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_CO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_CO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_CQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_C_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D5Q;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_DMUX;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_DO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_DO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_DQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_D_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X144Y121_SR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_AMUX;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_AO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_AO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_AQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_A_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B5Q;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_BMUX;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_BO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_BO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_BQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_B_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C5Q;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_CLK;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_CMUX;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_CO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_CO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_CQ;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_C_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D1;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D2;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D3;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D4;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_DO5;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_DO6;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D_CY;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_D_XOR;
  wire [0:0] CLBLM_L_X92Y121_SLICE_X145Y121_SR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_AO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_AO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_AQ;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_A_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B5Q;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_BMUX;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_BO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_BO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_BQ;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_B_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C5Q;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_CLK;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_CMUX;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_CO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_CO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_CQ;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_C_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_DO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_DO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_D_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X144Y122_SR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_AO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_AO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_AQ;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_A_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B5Q;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_BMUX;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_BO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_BO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_BQ;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_B_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C5Q;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_CLK;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_CMUX;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_CO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_CO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_CQ;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_C_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D1;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D2;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D3;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D4;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_DO5;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_DO6;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D_CY;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_D_XOR;
  wire [0:0] CLBLM_L_X92Y122_SLICE_X145Y122_SR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A5Q;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_AMUX;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_AO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_AO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_AQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_A_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_BO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_BO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_BQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_B_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_CLK;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_CO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_CO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_CQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_C_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D5Q;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_DMUX;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_DO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_DO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_DQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_D_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X144Y123_SR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A5Q;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_AMUX;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_AO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_AO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_AQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_A_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B5Q;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_BMUX;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_BO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_BO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_BQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_BX;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_B_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_CLK;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_CO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_CO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_CQ;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_C_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D1;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D2;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D3;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D4;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_DMUX;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_DO5;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_DO6;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D_CY;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_D_XOR;
  wire [0:0] CLBLM_L_X92Y123_SLICE_X145Y123_SR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A5Q;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_AMUX;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_AO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_AO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_AQ;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_AX;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_A_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_BMUX;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_BO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_BO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_B_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C5Q;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_CLK;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_CMUX;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_CO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_CO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_CQ;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_C_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_DO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_DO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_D_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X144Y124_SR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A5Q;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_AMUX;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_AO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_AO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_AQ;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_A_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_BO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_BO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_B_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_CLK;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_CO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_CO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_C_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D1;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D2;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D3;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D4;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_DO5;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_DO6;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D_CY;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_D_XOR;
  wire [0:0] CLBLM_L_X92Y124_SLICE_X145Y124_SR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_AO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_A_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_BO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_B_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_CO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_CO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_C_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_DO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_DO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X144Y125_D_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A5Q;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AMUX;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AQ;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_AX;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_A_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_BMUX;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_BO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_BO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_B_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C5Q;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CLK;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CMUX;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_CQ;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_C_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D1;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D2;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D3;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D4;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_DO5;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_DO6;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D_CY;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_D_XOR;
  wire [0:0] CLBLM_L_X92Y125_SLICE_X145Y125_SR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_AO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_AO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_AQ;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_AX;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_A_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_BO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_BO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_B_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_CLK;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_CO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_CO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_C_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_DO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_DO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_D_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X144Y126_SR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_AMUX;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_AO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_AO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_A_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B5Q;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_BMUX;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_BO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_BO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_BQ;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_B_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C5Q;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_CLK;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_CMUX;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_CO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_CO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_CQ;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_C_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D1;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D2;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D3;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D4;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_DO5;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_DO6;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D_CY;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_D_XOR;
  wire [0:0] CLBLM_L_X92Y126_SLICE_X145Y126_SR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_AO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_AO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_A_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_BO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_BO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_B_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_CO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_CO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_C_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_DO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_DO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X144Y127_D_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_AO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_AO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_AQ;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_A_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B5Q;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_BMUX;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_BO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_BO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_BQ;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_B_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_CLK;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_CO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_CO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_C_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D1;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D2;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D3;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D4;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_DO5;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_DO6;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D_CY;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_D_XOR;
  wire [0:0] CLBLM_L_X92Y127_SLICE_X145Y127_SR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_AO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_AO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_A_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_BO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_BO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_B_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_CO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_CO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_C_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_DO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_DO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X144Y128_D_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A5Q;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_AMUX;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_AO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_AO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_AQ;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_AX;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_A_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_BMUX;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_BO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_BO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_B_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C5Q;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_CLK;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_CMUX;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_CO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_CO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_CQ;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_C_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D1;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D2;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D3;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D4;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_DO5;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_DO6;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D_CY;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_D_XOR;
  wire [0:0] CLBLM_L_X92Y128_SLICE_X145Y128_SR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_AO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_AO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_A_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_BO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_BO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_B_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_CO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_CO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_C_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_DO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_DO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X144Y129_D_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A5Q;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_AMUX;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_AO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_AO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_AQ;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_AX;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_A_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_BMUX;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_BO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_BO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_B_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C5Q;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_CLK;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_CMUX;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_CO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_CO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_CQ;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_C_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D1;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D2;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D3;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D4;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_DO5;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_DO6;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D_CY;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_D_XOR;
  wire [0:0] CLBLM_L_X92Y129_SLICE_X145Y129_SR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A5Q;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_AMUX;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_AO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_AO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_AQ;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_A_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B5Q;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_BMUX;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_BO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_BO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_BQ;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_B_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C5Q;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_CLK;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_CMUX;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_CO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_CO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_CQ;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_C_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_DO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_DO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_D_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X144Y131_SR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A5Q;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_AMUX;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_AO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_AO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_AQ;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_AX;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_A_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_BMUX;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_BO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_BO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_B_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_CLK;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_CO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_CO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_C_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D1;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D2;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D3;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D4;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_DO5;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_DO6;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D_CY;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_D_XOR;
  wire [0:0] CLBLM_L_X92Y131_SLICE_X145Y131_SR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_AO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_AO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_A_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_BO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_BO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_B_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_CO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_CO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_C_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_DO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_DO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X144Y132_D_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A5Q;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_AMUX;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_AO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_AO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_AQ;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_AX;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_A_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_BMUX;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_BO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_BO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_B_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C5Q;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_CLK;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_CMUX;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_CO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_CO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_CQ;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_C_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D1;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D2;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D3;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D4;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_DO5;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_DO6;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D_CY;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_D_XOR;
  wire [0:0] CLBLM_L_X92Y132_SLICE_X145Y132_SR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_AO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_AO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_A_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_BO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_BO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_B_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_CO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_CO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_C_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_DO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_DO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X148Y111_D_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A5Q;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_AMUX;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_AO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_AO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_AQ;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_A_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B5Q;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_BMUX;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_BO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_BO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_BQ;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_B_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_CLK;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_CMUX;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_CO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_CO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_C_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D1;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D2;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D3;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D4;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_DO5;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_DO6;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D_CY;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_D_XOR;
  wire [0:0] CLBLM_L_X94Y111_SLICE_X149Y111_SR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A5Q;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_AMUX;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_AO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_AO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_AQ;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_A_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B5Q;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_BMUX;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_BO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_BO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_BQ;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_B_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_CLK;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_CO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_CO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_C_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_DO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_DO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_D_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X148Y112_SR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A5Q;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_AMUX;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_AO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_AO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_AQ;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_A_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B5Q;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_BMUX;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_BO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_BO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_BQ;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_B_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_CLK;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_CMUX;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_CO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_CO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_C_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D1;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D2;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D3;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D4;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_DO5;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_DO6;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D_CY;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_D_XOR;
  wire [0:0] CLBLM_L_X94Y112_SLICE_X149Y112_SR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A5Q;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_AMUX;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_AO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_AO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_AQ;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_A_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B5Q;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_BMUX;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_BO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_BO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_BQ;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_B_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_CLK;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_CO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_CO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_C_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_DO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_DO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_D_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X148Y113_SR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A5Q;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_AMUX;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_AO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_AO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_AQ;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_A_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_BMUX;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_BO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_BO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_B_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_CLK;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_CO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_CO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_C_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D1;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D2;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D3;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D4;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_DO5;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_DO6;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D_CY;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_D_XOR;
  wire [0:0] CLBLM_L_X94Y113_SLICE_X149Y113_SR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A5Q;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_AMUX;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_AO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_AO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_AQ;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_A_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B5Q;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_BMUX;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_BO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_BO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_BQ;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_B_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_CLK;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_CO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_CO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_C_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_DO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_DO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_D_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X148Y114_SR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A5Q;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_AMUX;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_AO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_AO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_AQ;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_A_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B5Q;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_BMUX;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_BO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_BO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_BQ;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_B_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_CLK;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_CO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_CO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_C_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D1;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D2;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D3;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D4;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_DMUX;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_DO5;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_DO6;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D_CY;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_D_XOR;
  wire [0:0] CLBLM_L_X94Y114_SLICE_X149Y114_SR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A5Q;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_AMUX;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_AO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_AO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_AQ;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_A_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B5Q;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_BMUX;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_BO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_BO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_BQ;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_B_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C5Q;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_CLK;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_CMUX;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_CO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_CO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_CQ;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_C_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_DMUX;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_DO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_DO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_D_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X148Y115_SR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A5Q;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_AMUX;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_AO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_AO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_AQ;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_A_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B5Q;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_BMUX;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_BO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_BO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_BQ;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_B_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_CLK;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_CO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_CO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_C_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D1;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D2;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D3;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D4;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_DO5;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_DO6;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D_CY;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_D_XOR;
  wire [0:0] CLBLM_L_X94Y115_SLICE_X149Y115_SR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A5Q;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_AMUX;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_AO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_AO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_AQ;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_A_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B5Q;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_BMUX;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_BO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_BO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_BQ;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_B_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_CLK;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_CO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_CO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_C_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_DMUX;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_DO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_DO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_D_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X148Y116_SR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A5Q;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_AMUX;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_AO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_AO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_AQ;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_A_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B5Q;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_BMUX;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_BO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_BO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_BQ;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_B_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C5Q;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_CLK;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_CMUX;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_CO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_CO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_CQ;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_C_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D1;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D2;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D3;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D4;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_DO5;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_DO6;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D_CY;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_D_XOR;
  wire [0:0] CLBLM_L_X94Y116_SLICE_X149Y116_SR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A5Q;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_AMUX;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_AO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_AO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_AQ;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_A_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B5Q;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_BMUX;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_BO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_BO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_BQ;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_B_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_CLK;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_CO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_CO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_C_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_DO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_DO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_D_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X148Y117_SR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A5Q;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_AMUX;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_AO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_AO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_AQ;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_A_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B5Q;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_BMUX;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_BO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_BO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_BQ;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_B_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_CLK;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_CO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_CO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_C_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D1;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D2;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D3;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D4;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_DO5;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_DO6;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D_CY;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_D_XOR;
  wire [0:0] CLBLM_L_X94Y117_SLICE_X149Y117_SR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A5Q;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_AMUX;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_AO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_AO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_AQ;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_A_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_BO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_BO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_B_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_CLK;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_CO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_CO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_C_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_DO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_DO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_D_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X148Y118_SR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A5Q;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_AMUX;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_AO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_AO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_AQ;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_A_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_BO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_BO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_B_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_CLK;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_CO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_CO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_C_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D1;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D2;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D3;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D4;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_DO5;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_DO6;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D_CY;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_D_XOR;
  wire [0:0] CLBLM_L_X94Y118_SLICE_X149Y118_SR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A5Q;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_AMUX;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_AO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_AO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_AQ;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_A_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_BO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_BO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_B_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_CLK;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_CMUX;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_CO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_CO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_C_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_DO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_DO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_D_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X148Y119_SR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A5Q;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_AMUX;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_AO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_AO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_AQ;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_A_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B5Q;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_BMUX;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_BO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_BO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_BQ;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_B_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_CLK;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_CO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_CO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_C_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D1;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D2;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D3;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D4;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_DO5;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_DO6;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D_CY;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_D_XOR;
  wire [0:0] CLBLM_L_X94Y119_SLICE_X149Y119_SR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A5Q;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_AMUX;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_AO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_AO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_AQ;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_A_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B5Q;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_BMUX;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_BO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_BO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_BQ;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_B_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C5Q;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_CLK;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_CMUX;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_CO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_CO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_CQ;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_C_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_DO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_DO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_D_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X148Y120_SR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A5Q;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_AMUX;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_AO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_AO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_AQ;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_A_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B5Q;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_BMUX;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_BO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_BO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_BQ;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_B_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_CLK;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_CMUX;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_CO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_CO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_C_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D1;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D2;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D3;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D4;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_DO5;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_DO6;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D_CY;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_D_XOR;
  wire [0:0] CLBLM_L_X94Y120_SLICE_X149Y120_SR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A5Q;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_AMUX;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_AO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_AO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_AQ;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_AX;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_A_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_BMUX;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_BO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_BO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_B_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C5Q;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_CLK;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_CMUX;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_CO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_CO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_CQ;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_C_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_DO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_DO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_D_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X148Y121_SR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A5Q;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_AMUX;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_AO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_AO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_AQ;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_A_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_BO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_BO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_B_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_CLK;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_CO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_CO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_C_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D1;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D2;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D3;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D4;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_DO5;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_DO6;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D_CY;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_D_XOR;
  wire [0:0] CLBLM_L_X94Y121_SLICE_X149Y121_SR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_AO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_A_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_BO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_B_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_CO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_CO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_C_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_DO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_DO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X148Y122_D_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A5Q;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_AMUX;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_AO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_AO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_AQ;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_A_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B5Q;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_BMUX;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_BO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_BO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_BQ;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_B_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_CLK;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_CO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_CO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_C_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D1;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D2;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D3;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D4;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_DO5;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_DO6;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D_CY;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_D_XOR;
  wire [0:0] CLBLM_L_X94Y122_SLICE_X149Y122_SR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A5Q;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_AMUX;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_AO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_AO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_AQ;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_AX;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_A_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_BMUX;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_BO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_BO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_B_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C5Q;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_CLK;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_CMUX;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_CO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_CO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_CQ;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_C_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_DO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_DO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_D_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X148Y123_SR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_AO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_AO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_A_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_BO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_BO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_B_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_CO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_CO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_C_XOR;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D1;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D2;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D3;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D4;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_DO5;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_DO6;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D_CY;
  wire [0:0] CLBLM_L_X94Y123_SLICE_X149Y123_D_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A5Q;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_AMUX;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_AO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_AO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_AQ;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_A_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B5Q;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_BMUX;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_BO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_BO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_BQ;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_B_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C5Q;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_CLK;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_CMUX;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_CO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_CO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_CQ;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_C_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_DO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_DO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_D_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X148Y124_SR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A5Q;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_AMUX;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_AO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_AO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_AQ;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_A_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_BO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_BO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_B_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_CLK;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_CO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_CO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_C_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D1;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D2;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D3;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D4;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_DO5;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_DO6;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D_CY;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_D_XOR;
  wire [0:0] CLBLM_L_X94Y124_SLICE_X149Y124_SR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A5Q;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_AMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_AO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_AO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_AQ;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_A_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B5Q;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_BMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_BO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_BO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_BQ;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_B_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_CLK;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_CMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_CO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_CO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_C_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_DO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_DO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_D_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X148Y125_SR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A5Q;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_AMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_AO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_AO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_AQ;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_AX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_A_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_BMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_BO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_BO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_B_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C5Q;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_CLK;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_CMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_CO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_CO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_CQ;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_C_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D1;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D2;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D3;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D4;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D5Q;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_DMUX;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_DO5;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_DO6;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_DQ;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D_CY;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_D_XOR;
  wire [0:0] CLBLM_L_X94Y125_SLICE_X149Y125_SR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_AO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_AO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_A_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_BO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_BO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_B_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_CO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_CO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_C_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_DO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_DO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X148Y126_D_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_AO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_AO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_A_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_BO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_BO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_B_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_CO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_CO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_C_XOR;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D1;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D2;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D3;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D4;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_DO5;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_DO6;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D_CY;
  wire [0:0] CLBLM_L_X94Y126_SLICE_X149Y126_D_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_AO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_AO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_A_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_BO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_BO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_B_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_CO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_CO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_C_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_DO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_DO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X148Y127_D_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A5Q;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_AMUX;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_AO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_AO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_AQ;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_A_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B5Q;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_BMUX;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_BO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_BO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_BQ;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_BX;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_B_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_CLK;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_CMUX;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_CO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_CO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_C_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D1;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D2;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D3;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D4;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_DO5;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_DO6;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D_CY;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_D_XOR;
  wire [0:0] CLBLM_L_X94Y127_SLICE_X149Y127_SR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_AO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_AO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_A_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_BO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_BO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_B_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_CO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_CO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_C_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_DO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_DO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X148Y128_D_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A5Q;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_AMUX;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_AO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_AO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_AQ;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_AX;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_A_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_BMUX;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_BO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_BO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_B_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C5Q;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_CLK;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_CMUX;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_CO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_CO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_CQ;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_C_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D1;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D2;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D3;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D4;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_DO5;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_DO6;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D_CY;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_D_XOR;
  wire [0:0] CLBLM_L_X94Y128_SLICE_X149Y128_SR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_AO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_AO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_AQ;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_A_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B5Q;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_BMUX;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_BO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_BO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_BQ;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_B_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_CLK;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_CO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_CO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_C_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_DO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_DO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_D_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X148Y129_SR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_AO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_AO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_A_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_BO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_BO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_B_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_CO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_CO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_C_XOR;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D1;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D2;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D3;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D4;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_DO5;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_DO6;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D_CY;
  wire [0:0] CLBLM_L_X94Y129_SLICE_X149Y129_D_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_AO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_AO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_AQ;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_A_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_BO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_BO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_B_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_CLK;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_CO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_CO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_C_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_DO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_DO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_D_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X148Y130_SR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A5Q;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_AMUX;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_AO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_AO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_AQ;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_A_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_BO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_BO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_B_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_CLK;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_CO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_CO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_C_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D1;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D2;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D3;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D4;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_DO5;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_DO6;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D_CY;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_D_XOR;
  wire [0:0] CLBLM_L_X94Y130_SLICE_X149Y130_SR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_AO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_AO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_A_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_BO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_BO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_B_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_CO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_CO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_C_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_DO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_DO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X148Y132_D_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_AMUX;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_AO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_AO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_A_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_BO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_BO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_B_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_CO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_CO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_C_XOR;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D1;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D2;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D3;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D4;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_DO5;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_DO6;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D_CY;
  wire [0:0] CLBLM_L_X94Y132_SLICE_X149Y132_D_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A5Q;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_AMUX;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_AO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_AO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_AQ;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_A_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_BO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_BO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_B_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_CLK;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_CO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_CO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_C_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_DO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_DO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_D_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X154Y110_SR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_AO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_AO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_A_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_BO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_BO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_B_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_CO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_CO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_C_XOR;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D1;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D2;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D3;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D4;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_DO5;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_DO6;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D_CY;
  wire [0:0] CLBLM_L_X98Y110_SLICE_X155Y110_D_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A5Q;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_AMUX;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_AO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_AO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_AQ;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_A_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B5Q;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_BMUX;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_BO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_BO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_BQ;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_B_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_CLK;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_CO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_CO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_C_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_DO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_DO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_D_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X154Y111_SR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A5Q;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_AMUX;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_AO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_AO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_AQ;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_A_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B5Q;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_BMUX;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_BO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_BO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_BQ;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_B_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C5Q;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_CLK;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_CMUX;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_CO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_CO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_CQ;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_C_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D1;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D2;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D3;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D4;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_DMUX;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_DO5;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_DO6;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D_CY;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_D_XOR;
  wire [0:0] CLBLM_L_X98Y111_SLICE_X155Y111_SR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A5Q;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_AMUX;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_AO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_AO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_AQ;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_A_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B5Q;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_BMUX;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_BO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_BO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_BQ;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_B_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_CLK;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_CMUX;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_CO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_CO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_C_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_DO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_DO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_D_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X154Y112_SR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A5Q;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_AMUX;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_AO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_AO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_AQ;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_A_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_BO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_BO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_B_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_CLK;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_CO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_CO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_C_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D1;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D2;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D3;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D4;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_DO5;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_DO6;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D_CY;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_D_XOR;
  wire [0:0] CLBLM_L_X98Y112_SLICE_X155Y112_SR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A5Q;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_AMUX;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_AO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_AO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_AQ;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_A_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_BO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_BO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_B_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_CLK;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_CO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_CO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_C_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_DO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_DO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_D_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X154Y113_SR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_AO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_AO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_A_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_BO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_BO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_B_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_CO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_CO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_C_XOR;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D1;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D2;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D3;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D4;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_DO5;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_DO6;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D_CY;
  wire [0:0] CLBLM_L_X98Y113_SLICE_X155Y113_D_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A5Q;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_AMUX;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_AO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_AO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_AQ;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_A_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B5Q;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_BMUX;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_BO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_BO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_BQ;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_B_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C5Q;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_CLK;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_CMUX;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_CO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_CO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_CQ;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_C_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_DO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_DO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_D_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X154Y114_SR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_AO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_AO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_A_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_BO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_BO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_B_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_CO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_CO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_C_XOR;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D1;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D2;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D3;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D4;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_DO5;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_DO6;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D_CY;
  wire [0:0] CLBLM_L_X98Y114_SLICE_X155Y114_D_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A5Q;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_AMUX;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_AO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_AO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_AQ;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_A_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B5Q;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_BMUX;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_BO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_BO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_BQ;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_B_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_CLK;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_CO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_CO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_C_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_DO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_DO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_D_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X154Y115_SR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A5Q;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_AMUX;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_AO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_AO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_AQ;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_A_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B5Q;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_BMUX;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_BO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_BO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_BQ;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_B_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C5Q;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_CLK;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_CMUX;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_CO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_CO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_CQ;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_C_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D1;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D2;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D3;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D4;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_DO5;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_DO6;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D_CY;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_D_XOR;
  wire [0:0] CLBLM_L_X98Y115_SLICE_X155Y115_SR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_AO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_AO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_A_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_BO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_BO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_B_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_CO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_CO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_C_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_DO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_DO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X154Y116_D_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A5Q;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_AMUX;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_AO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_AO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_AQ;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_A_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B5Q;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_BMUX;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_BO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_BO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_BQ;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_B_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_CLK;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_CO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_CO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_C_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D1;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D2;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D3;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D4;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_DO5;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_DO6;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D_CY;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_D_XOR;
  wire [0:0] CLBLM_L_X98Y116_SLICE_X155Y116_SR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_AO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_AO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_A_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_BO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_BO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_B_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_CO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_CO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_C_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_DO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_DO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X154Y117_D_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A5Q;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_AMUX;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_AO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_AO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_AQ;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_A_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B5Q;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_BMUX;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_BO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_BO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_BQ;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_B_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_CLK;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_CO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_CO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_C_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D1;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D2;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D3;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D4;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_DO5;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_DO6;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D_CY;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_D_XOR;
  wire [0:0] CLBLM_L_X98Y117_SLICE_X155Y117_SR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A5Q;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_AMUX;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_AO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_AO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_AQ;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_A_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B5Q;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_BMUX;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_BO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_BO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_BQ;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_BX;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_B_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_CLK;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_CMUX;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_CO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_CO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_C_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_DO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_DO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_D_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X154Y119_SR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_AO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_AO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_AQ;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_A_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B5Q;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_BMUX;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_BO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_BO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_BQ;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_B_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C5Q;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_CLK;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_CMUX;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_CO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_CO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_CQ;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_C_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D1;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D2;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D3;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D4;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_DO5;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_DO6;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D_CY;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_D_XOR;
  wire [0:0] CLBLM_L_X98Y119_SLICE_X155Y119_SR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A5Q;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_AMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_AO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_AO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_AQ;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_AX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_A_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_BMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_BO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_BO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_B_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C5Q;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_CLK;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_CMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_CO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_CO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_CQ;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_C_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_DMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_DO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_DO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_D_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X154Y120_SR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A5Q;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_AMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_AO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_AO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_AQ;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_A_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B5Q;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_BMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_BO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_BO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_BQ;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_B_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_CLK;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_CO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_CO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_C_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D1;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D2;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D3;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D4;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_DMUX;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_DO5;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_DO6;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D_CY;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_D_XOR;
  wire [0:0] CLBLM_L_X98Y120_SLICE_X155Y120_SR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A5Q;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_AMUX;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_AO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_AO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_AQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_A_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_BO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_BO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_BQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_B_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_CLK;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_CO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_CO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_CQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_C_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D5Q;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_DMUX;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_DO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_DO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_DQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_D_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X154Y121_SR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_AO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_AO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_AQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_A_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B5Q;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_BMUX;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_BO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_BO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_BQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_B_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C5Q;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_CLK;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_CMUX;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_CO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_CO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_CQ;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_C_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D1;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D2;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D3;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D4;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_DO5;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_DO6;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D_CY;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_D_XOR;
  wire [0:0] CLBLM_L_X98Y121_SLICE_X155Y121_SR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A5Q;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_AMUX;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_AO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_AO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_AQ;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_A_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B5Q;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_BMUX;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_BO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_BO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_BQ;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_B_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_CLK;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_CO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_CO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_C_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_DO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_DO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_D_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X154Y122_SR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A5Q;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_AMUX;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_AO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_AO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_AQ;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_A_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B5Q;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_BMUX;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_BO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_BO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_BQ;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_B_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_CLK;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_CO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_CO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_C_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D1;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D2;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D3;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D4;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_DO5;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_DO6;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D_CY;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_D_XOR;
  wire [0:0] CLBLM_L_X98Y122_SLICE_X155Y122_SR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A5Q;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_AMUX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_AO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_AO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_AQ;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_AX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_A_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_BMUX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_BO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_BO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_B_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C5Q;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_CLK;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_CMUX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_CO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_CO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_CQ;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_C_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_DO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_DO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_D_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X154Y123_SR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A5Q;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_AMUX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_AO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_AO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_AQ;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_AX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_A_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_BMUX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_BO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_BO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_B_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C5Q;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_CLK;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_CMUX;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_CO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_CO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_CQ;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_C_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D1;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D2;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D3;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D4;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_DO5;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_DO6;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D_CY;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_D_XOR;
  wire [0:0] CLBLM_L_X98Y123_SLICE_X155Y123_SR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A5Q;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_AMUX;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_AO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_AO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_AQ;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_A_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B5Q;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_BMUX;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_BO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_BO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_BQ;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_B_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_CLK;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_CO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_CO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_C_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_DO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_DO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_D_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X154Y124_SR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_AO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_AO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_A_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_BO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_BO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_B_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_CO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_CO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_C_XOR;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D1;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D2;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D3;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D4;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_DO5;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_DO6;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D_CY;
  wire [0:0] CLBLM_L_X98Y124_SLICE_X155Y124_D_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A5Q;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_AMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_AO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_AO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_AQ;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_A_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B5Q;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_BMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_BO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_BO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_BQ;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_B_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C5Q;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_CLK;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_CMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_CO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_CO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_CQ;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_C_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D5Q;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_DMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_DO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_DO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_DQ;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_D_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X154Y125_SR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A5Q;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_AMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_AO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_AO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_AQ;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_AX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_A_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_BMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_BO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_BO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_B_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C5Q;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_CLK;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_CMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_CO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_CO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_CQ;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_C_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D1;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D2;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D3;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D4;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_DMUX;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_DO5;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_DO6;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D_CY;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_D_XOR;
  wire [0:0] CLBLM_L_X98Y125_SLICE_X155Y125_SR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A5Q;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_AMUX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_AO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_AO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_AQ;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_A_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B5Q;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_BMUX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_BO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_BO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_BQ;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_B_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_CLK;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_CMUX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_CO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_CO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_C_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_DO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_DO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_D_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X154Y126_SR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A5Q;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_AMUX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_AO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_AO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_AQ;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_AX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_A_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_BMUX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_BO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_BO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_B_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C5Q;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_CLK;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_CMUX;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_CO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_CO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_CQ;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_C_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D1;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D2;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D3;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D4;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_DO5;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_DO6;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D_CY;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_D_XOR;
  wire [0:0] CLBLM_L_X98Y126_SLICE_X155Y126_SR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A5Q;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_AMUX;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_AO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_AO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_AQ;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_A_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B5Q;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_BMUX;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_BO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_BO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_BQ;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_B_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_CLK;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_CMUX;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_CO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_CO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_C_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_DO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_DO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_D_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X154Y127_SR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A5Q;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_AMUX;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_AO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_AO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_AQ;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_A_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B5Q;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_BMUX;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_BO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_BO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_BQ;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_B_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_CLK;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_CO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_CO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_C_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D1;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D2;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D3;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D4;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_DO5;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_DO6;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D_CY;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_D_XOR;
  wire [0:0] CLBLM_L_X98Y127_SLICE_X155Y127_SR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A5Q;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_AMUX;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_AO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_AO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_AQ;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_A_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B5Q;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_BMUX;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_BO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_BO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_BQ;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_B_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C5Q;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_CLK;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_CMUX;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_CO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_CO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_CQ;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_C_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_DO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_DO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_D_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X154Y128_SR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_AO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_AO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_A_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_BO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_BO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_B_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_CO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_CO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_C_XOR;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D1;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D2;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D3;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D4;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_DO5;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_DO6;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D_CY;
  wire [0:0] CLBLM_L_X98Y128_SLICE_X155Y128_D_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_AMUX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_AO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_AO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_AQ;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_AX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_A_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B5Q;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_BMUX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_BO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_BO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_BQ;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_B_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_CLK;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_CO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_CO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_CQ;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_CX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_C_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_DO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_DO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_D_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X154Y129_SR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A5Q;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_AMUX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_AO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_AO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_AQ;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_A_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_BMUX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_BO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_BO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_B_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C5Q;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_CLK;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_CMUX;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_CO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_CO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_CQ;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_C_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D1;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D2;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D3;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D4;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_DO5;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_DO6;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D_CY;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_D_XOR;
  wire [0:0] CLBLM_L_X98Y129_SLICE_X155Y129_SR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A5Q;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_AMUX;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_AO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_AO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_AQ;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_AX;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_A_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_BMUX;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_BO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_BO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_B_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C5Q;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_CLK;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_CMUX;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_CO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_CO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_CQ;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_C_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_DO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_DO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_D_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X154Y130_SR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A5Q;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_AMUX;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_AO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_AO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_AQ;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_A_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_BO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_BO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_BQ;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_B_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_CLK;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_CO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_CO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_CQ;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_C_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D1;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D2;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D3;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D4;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D5Q;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_DMUX;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_DO5;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_DO6;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_DQ;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D_CY;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_D_XOR;
  wire [0:0] CLBLM_L_X98Y130_SLICE_X155Y130_SR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A5Q;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AQ;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_BMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_BO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_BO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C5Q;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CLK;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CQ;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_DO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_DO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_SR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A5Q;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_AMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_AO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_AO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_AQ;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B5Q;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BQ;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_CLK;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_CMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_CO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_CO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D5Q;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_DMUX;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_DO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_DO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_DQ;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_SR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A5Q;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AMUX;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AQ;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AX;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_BMUX;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_BO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_BO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C5Q;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CLK;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CMUX;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CQ;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_DO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_DO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_SR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_AO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_AO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_AQ;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_BO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_BO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_BQ;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C5Q;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CLK;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CMUX;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CQ;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_DO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_DO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_SR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A5Q;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_AMUX;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_AO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_AO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_AQ;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_A_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B5Q;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_BMUX;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_BO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_BO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_BQ;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_B_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_CLK;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_CO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_CO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_C_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_DO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_DO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_D_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X154Y133_SR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A5Q;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_AMUX;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_AO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_AO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_AQ;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_A_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_BO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_BO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_BQ;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_B_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_CLK;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_CO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_CO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_C_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D1;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D2;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D3;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D4;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_DO5;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_DO6;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D_CY;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_D_XOR;
  wire [0:0] CLBLM_L_X98Y133_SLICE_X155Y133_SR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A5Q;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_AMUX;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_AO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_AO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_AQ;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_AX;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_A_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_BMUX;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_BO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_BO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_B_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C5Q;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_CLK;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_CMUX;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_CO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_CO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_CQ;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_C_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_DO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_DO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_D_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X154Y134_SR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_AO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_AO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_A_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_BO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_BO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_B_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_CO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_CO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_C_XOR;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D1;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D2;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D3;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D4;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_DO5;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_DO6;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D_CY;
  wire [0:0] CLBLM_L_X98Y134_SLICE_X155Y134_D_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A5Q;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_AMUX;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_AO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_AO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_AQ;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_A_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B5Q;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_BMUX;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_BO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_BO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_BQ;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_B_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_CLK;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_CO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_CO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_C_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_DO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_DO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_D_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X158Y110_SR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_AO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_AO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_A_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_BO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_BO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_B_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_CO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_CO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_C_XOR;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D1;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D2;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D3;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D4;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_DO5;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_DO6;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D_CY;
  wire [0:0] CLBLM_R_X101Y110_SLICE_X159Y110_D_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A5Q;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_AMUX;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_AO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_AO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_AQ;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_A_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B5Q;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_BMUX;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_BO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_BO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_BQ;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_B_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_CLK;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_CMUX;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_CO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_CO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_C_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_DO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_DO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_D_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X158Y111_SR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A5Q;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_AMUX;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_AO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_AO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_AQ;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_A_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B5Q;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_BMUX;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_BO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_BO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_BQ;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_B_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_CLK;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_CO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_CO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_C_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D1;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D2;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D3;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D4;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_DO5;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_DO6;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D_CY;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_D_XOR;
  wire [0:0] CLBLM_R_X101Y111_SLICE_X159Y111_SR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A5Q;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_AMUX;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_AO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_AO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_AQ;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_A_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B5Q;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_BMUX;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_BO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_BO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_BQ;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_B_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_CLK;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_CO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_CO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_C_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_DO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_DO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_D_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X158Y112_SR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A5Q;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_AMUX;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_AO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_AO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_AQ;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_A_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B5Q;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_BMUX;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_BO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_BO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_BQ;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_B_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C5Q;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_CLK;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_CMUX;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_CO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_CO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_CQ;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_C_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D1;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D2;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D3;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D4;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_DO5;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_DO6;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D_CY;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_D_XOR;
  wire [0:0] CLBLM_R_X101Y112_SLICE_X159Y112_SR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A5Q;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_AMUX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_AO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_AO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_AQ;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_A_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B5Q;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_BMUX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_BO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_BO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_BQ;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_B_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_CLK;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_CO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_CO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_C_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_DO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_DO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_D_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X158Y113_SR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_AMUX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_AO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_AO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_AQ;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_AX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_A_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_BMUX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_BO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_BO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_BQ;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_BX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_B_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C5Q;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_CLK;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_CMUX;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_CO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_CO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_CQ;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_C_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D1;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D2;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D3;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D4;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_DO5;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_DO6;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D_CY;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_D_XOR;
  wire [0:0] CLBLM_R_X101Y113_SLICE_X159Y113_SR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A5Q;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_AMUX;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_AO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_AO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_AQ;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_A_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B5Q;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_BMUX;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_BO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_BO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_BQ;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_B_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_CLK;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_CMUX;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_CO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_CO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_C_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_DO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_DO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_D_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X158Y114_SR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_AO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_AO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_A_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_BO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_BO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_B_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_CO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_CO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_C_XOR;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D1;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D2;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D3;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D4;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_DO5;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_DO6;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D_CY;
  wire [0:0] CLBLM_R_X101Y114_SLICE_X159Y114_D_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A5Q;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_AMUX;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_AO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_AO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_AQ;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_A_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B5Q;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_BMUX;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_BO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_BO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_BQ;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_B_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_CLK;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_CO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_CO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_C_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_DO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_DO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_D_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X158Y115_SR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_AO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_AO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_A_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_BO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_BO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_B_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_CO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_CO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_C_XOR;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D1;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D2;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D3;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D4;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_DO5;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_DO6;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D_CY;
  wire [0:0] CLBLM_R_X101Y115_SLICE_X159Y115_D_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A5Q;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_AMUX;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_AO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_AO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_AQ;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B5Q;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_BMUX;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_BO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_BO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_BQ;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_CLK;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_CMUX;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_CO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_CO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_DO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_DO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_SR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_AMUX;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_AO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_BMUX;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_BO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C5Q;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CLK;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CMUX;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CQ;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_DO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_DO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_SR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_AO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_AO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_AQ;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B5Q;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_BMUX;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_BO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_BO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_BQ;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_CLK;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_CMUX;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_CO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_CO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_DO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_DO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_SR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_AMUX;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_AO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_AO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_AQ;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B5Q;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_BMUX;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_BO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_BO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_BQ;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_CLK;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_CO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_CO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_CQ;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_DO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_DO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_SR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A5Q;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_AMUX;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_AO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_AQ;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B5Q;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_BMUX;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_BO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_BQ;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_CLK;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_CO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_CQ;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_DO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_SR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A5Q;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_AMUX;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_AO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_AO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_AQ;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B5Q;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_BMUX;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_BO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_BO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_BQ;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CLK;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CMUX;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CQ;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CX;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_DO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_DO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_SR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A5Q;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_AMUX;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_AO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_AQ;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_BO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_BQ;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_CLK;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_CO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_CQ;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_DO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_SR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A5Q;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_AMUX;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_AO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_AO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_AQ;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B5Q;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_BMUX;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_BO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_BO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_BQ;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_CLK;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_CO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_DO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_DO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_SR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A5Q;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_AMUX;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_AO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_AO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_AQ;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_AX;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_A_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_BMUX;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_BO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_BO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_B_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C5Q;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_CLK;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_CMUX;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_CO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_CO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_CQ;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_C_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_DMUX;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_DO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_DO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_D_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X158Y120_SR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_AO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_AO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_AQ;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_A_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B5Q;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_BMUX;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_BO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_BO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_BQ;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_B_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_CLK;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_CO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_CO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_C_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D1;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D2;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D3;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D4;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_DO5;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_DO6;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D_CY;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_D_XOR;
  wire [0:0] CLBLM_R_X101Y120_SLICE_X159Y120_SR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A5Q;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_AMUX;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_AO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_AO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_AQ;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_A_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_BO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_BO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_B_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_CLK;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_CO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_CO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_C_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_DO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_DO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_D_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X158Y121_SR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A5Q;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_AMUX;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_AO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_AO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_AQ;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_A_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B5Q;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_BMUX;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_BO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_BO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_BQ;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_B_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C5Q;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_CLK;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_CMUX;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_CO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_CO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_CQ;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_C_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D1;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D2;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D3;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D4;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_DMUX;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_DO5;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_DO6;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D_CY;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_D_XOR;
  wire [0:0] CLBLM_R_X101Y121_SLICE_X159Y121_SR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A5Q;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_AMUX;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_AO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_AO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_AQ;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_A_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B5Q;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_BMUX;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_BO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_BO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_BQ;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_B_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_CLK;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_CO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_CO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_C_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_DMUX;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_DO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_DO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_D_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X158Y122_SR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A5Q;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_AMUX;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_AO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_AO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_AQ;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_A_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B5Q;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_BMUX;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_BO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_BO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_BQ;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_B_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_CLK;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_CO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_CO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_C_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D1;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D2;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D3;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D4;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_DO5;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_DO6;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D_CY;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_D_XOR;
  wire [0:0] CLBLM_R_X101Y122_SLICE_X159Y122_SR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A5Q;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AQ;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B5Q;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BQ;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CLK;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_SR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A5Q;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AQ;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BQ;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C5Q;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CLK;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CQ;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_DO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_DO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_SR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A5Q;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_AMUX;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_AO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_AQ;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_A_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B5Q;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_BMUX;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_BO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_BQ;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_B_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_CLK;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_CMUX;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_CO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_C_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_DO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_D_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X158Y124_SR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A5Q;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_AMUX;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_AO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_AO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_AQ;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_A_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_BO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_BO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_B_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_CLK;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_CO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_CO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_C_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D1;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D2;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D3;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D4;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_DO5;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_DO6;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D_CY;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_D_XOR;
  wire [0:0] CLBLM_R_X101Y124_SLICE_X159Y124_SR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_AO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_AO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_AQ;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_A_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B5Q;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_BMUX;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_BO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_BO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_BQ;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_B_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_CLK;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_CO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_CO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_C_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_DO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_DO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_D_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X158Y125_SR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_AO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_AO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_A_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_BO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_BO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_B_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_CO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_CO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_C_XOR;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D1;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D2;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D3;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D4;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_DO5;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_DO6;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D_CY;
  wire [0:0] CLBLM_R_X101Y125_SLICE_X159Y125_D_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A5Q;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_AMUX;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_AO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_AO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_AQ;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_A_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_BO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_BO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_B_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_CLK;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_CO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_CO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_C_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_DO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_DO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_D_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X158Y126_SR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A5Q;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_AMUX;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_AO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_AO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_AQ;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_A_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_BO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_BO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_B_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_CLK;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_CO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_CO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_C_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D1;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D2;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D3;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D4;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_DO5;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_DO6;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D_CY;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_D_XOR;
  wire [0:0] CLBLM_R_X101Y126_SLICE_X159Y126_SR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_AO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_AO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_A_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_BO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_BO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_B_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_CO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_CO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_C_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_DO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_DO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X158Y127_D_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A5Q;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_AMUX;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_AO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_AO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_AQ;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_A_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_BO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_BO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_B_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_CLK;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_CO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_CO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_C_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D1;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D2;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D3;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D4;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_DO5;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_DO6;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D_CY;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_D_XOR;
  wire [0:0] CLBLM_R_X101Y127_SLICE_X159Y127_SR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A5Q;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_AMUX;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_AO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_AO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_AQ;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_A_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_BO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_BO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_B_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_CLK;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_CO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_CO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_C_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_DO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_DO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_D_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X158Y128_SR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_AO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_AO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_A_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_BO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_BO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_B_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_CO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_CO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_C_XOR;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D1;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D2;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D3;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D4;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_DO5;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_DO6;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D_CY;
  wire [0:0] CLBLM_R_X101Y128_SLICE_X159Y128_D_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A5Q;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_AMUX;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_AO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_AO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_AQ;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_A_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B5Q;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_BMUX;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_BO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_BO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_BQ;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_B_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_CLK;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_CO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_CO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_C_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_DO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_DO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_D_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X158Y129_SR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_AO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_AO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_AQ;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_A_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_BO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_BO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_B_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_CLK;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_CO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_CO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_C_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D1;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D2;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D3;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D4;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_DO5;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_DO6;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D_CY;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_D_XOR;
  wire [0:0] CLBLM_R_X101Y129_SLICE_X159Y129_SR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A5Q;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_AMUX;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_AO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_AO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_AQ;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_A_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_BO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_BO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_BQ;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_B_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C5Q;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_CLK;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_CMUX;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_CO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_CO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_CQ;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_C_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_DO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_DO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_D_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X158Y130_SR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_AO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_AO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_AQ;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_A_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B5Q;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_BMUX;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_BO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_BO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_BQ;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_B_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_CLK;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_CMUX;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_CO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_CO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_C_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D1;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D2;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D3;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D4;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_DO5;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_DO6;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D_CY;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_D_XOR;
  wire [0:0] CLBLM_R_X101Y130_SLICE_X159Y130_SR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_AO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_AO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_AQ;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_A_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B5Q;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_BMUX;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_BO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_BO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_BQ;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_B_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_CLK;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_CMUX;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_CO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_CO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_C_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_DO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_DO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_D_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X158Y131_SR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A5Q;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_AMUX;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_AO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_AO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_AQ;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_A_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B5Q;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_BMUX;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_BO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_BO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_BQ;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_B_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C5Q;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_CLK;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_CMUX;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_CO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_CO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_CQ;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_C_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D1;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D2;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D3;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D4;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D5Q;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_DMUX;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_DO5;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_DO6;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_DQ;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D_CY;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_D_XOR;
  wire [0:0] CLBLM_R_X101Y131_SLICE_X159Y131_SR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A5Q;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_AMUX;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_AO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_AO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_AQ;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_A_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_BO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_BO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_B_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_CLK;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_CO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_CO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_C_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_DO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_DO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_D_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X158Y132_SR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_AO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_AO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_AQ;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_A_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B5Q;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_BMUX;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_BO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_BO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_BQ;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_B_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_CLK;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_CMUX;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_CO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_CO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_C_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D1;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D2;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D3;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D4;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_DO5;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_DO6;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D_CY;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_D_XOR;
  wire [0:0] CLBLM_R_X101Y132_SLICE_X159Y132_SR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_AO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_AO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_AQ;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_A_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B5Q;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_BMUX;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_BO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_BO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_BQ;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_B_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_CLK;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_CO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_CO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_C_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_DO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_DO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_D_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X158Y133_SR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A5Q;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_AMUX;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_AO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_AO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_AQ;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_A_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_BO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_BO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_B_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_CLK;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_CO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_CO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_C_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D1;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D2;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D3;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D4;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_DO5;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_DO6;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D_CY;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_D_XOR;
  wire [0:0] CLBLM_R_X101Y133_SLICE_X159Y133_SR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A5Q;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_AMUX;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_AO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_AO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_AQ;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_A_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_BO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_BO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_B_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_CLK;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_CO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_CO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_C_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_DO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_DO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_D_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X158Y134_SR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_AO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_AO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_AQ;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_A_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_BO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_BO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_BQ;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_B_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C5Q;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_CLK;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_CMUX;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_CO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_CO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_CQ;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_C_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D1;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D2;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D3;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D4;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_DO5;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_DO6;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D_CY;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_D_XOR;
  wire [0:0] CLBLM_R_X101Y134_SLICE_X159Y134_SR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A5Q;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_AMUX;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_AO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_AO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_AQ;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_A_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_BO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_BO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_B_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_CLK;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_CO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_CO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_C_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_DO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_DO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_D_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X158Y135_SR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A5Q;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_AMUX;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_AO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_AO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_AQ;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_A_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B5Q;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_BMUX;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_BO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_BO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_BQ;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_B_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C5Q;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_CLK;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_CMUX;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_CO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_CO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_CQ;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_C_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D1;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D2;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D3;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D4;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D5Q;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_DMUX;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_DO5;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_DO6;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_DQ;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D_CY;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_D_XOR;
  wire [0:0] CLBLM_R_X101Y135_SLICE_X159Y135_SR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A5Q;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_AMUX;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_AO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_AO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_AQ;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_A_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_BO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_BO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_B_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_CLK;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_CO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_CO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_C_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_DO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_DO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_D_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X158Y136_SR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_AO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_AO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_AQ;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_A_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B5Q;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_BMUX;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_BO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_BO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_BQ;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_B_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_CLK;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_CO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_CO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_C_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D1;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D2;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D3;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D4;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_DO5;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_DO6;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D_CY;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_D_XOR;
  wire [0:0] CLBLM_R_X101Y136_SLICE_X159Y136_SR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AMUX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BMUX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CLK;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CMUX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_DO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_DO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_SR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_AO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_AO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_BO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_BO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_DO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_DO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AMUX;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B5Q;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_BMUX;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_BO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_BO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_BQ;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C5Q;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CLK;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CMUX;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CQ;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_DO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_DO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_SR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A5Q;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_AMUX;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_AO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_AO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_AQ;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_BO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_BO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_BQ;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_BX;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_CLK;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_CO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_CO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_DO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_DO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_SR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AMUX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BMUX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CLK;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_DO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_DO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_SR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BMUX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CLK;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_DO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_DO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_SR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CLK;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_DMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_DO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_SR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_AO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_AO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_CO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_DO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_DO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_AO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_AO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B5Q;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_BMUX;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_BO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_BQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_CLK;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_CO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_DO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_DO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_SR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_AO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_AO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_BO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_BO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_CO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_CO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_DO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_DO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AX;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_BO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_BO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_CLK;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_CO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_DO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_DO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_SR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_AO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_AO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_AQ;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B5Q;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_BMUX;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_BO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_BO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_BQ;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_CLK;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_CO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_DO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_DO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_SR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A5Q;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_AMUX;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_AO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_AO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_AQ;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_A_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B5Q;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_BMUX;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_BO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_BO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_BQ;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_B_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C5Q;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_CLK;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_CMUX;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_CO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_CO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_CQ;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_C_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_DO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_DO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_D_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X162Y120_SR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_AO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_AO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_AQ;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_A_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B5Q;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_BMUX;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_BO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_BO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_BQ;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_B_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_CLK;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_CO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_CO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_C_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D1;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D2;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D3;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D4;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_DO5;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_DO6;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D_CY;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_D_XOR;
  wire [0:0] CLBLM_R_X103Y120_SLICE_X163Y120_SR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_AO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_AO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_AQ;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_A_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B5Q;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_BMUX;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_BO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_BO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_BQ;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_B_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_CLK;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_CO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_CO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_C_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_DO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_DO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_D_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X162Y121_SR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A5Q;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_AMUX;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_AO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_AO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_AQ;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_A_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B5Q;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_BMUX;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_BO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_BO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_BQ;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_B_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C5Q;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_CLK;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_CMUX;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_CO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_CO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_CQ;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_C_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D1;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D2;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D3;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D4;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_DO5;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_DO6;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D_CY;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_D_XOR;
  wire [0:0] CLBLM_R_X103Y121_SLICE_X163Y121_SR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A5Q;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AQ;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B5Q;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BQ;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CLK;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_SR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A5Q;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B5Q;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BQ;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C5Q;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CLK;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CQ;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_SR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A5Q;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_AMUX;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_AO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_AQ;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_BO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_BQ;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_CLK;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_CO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_CQ;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_DO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_SR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_AO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_AO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_AQ;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_BO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_BO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_CLK;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_CO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_CO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_DO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_DO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_SR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_AO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_AO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_AQ;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_A_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B5Q;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_BMUX;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_BO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_BO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_BQ;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_B_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_CLK;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_CO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_CO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_C_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_DMUX;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_DO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_DO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_D_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X162Y124_SR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_AO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_AO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_AQ;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_A_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B5Q;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_BMUX;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_BO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_BO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_BQ;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_B_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_CLK;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_CO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_CO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_C_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D1;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D2;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D3;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D4;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_DMUX;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_DO5;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_DO6;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D_CY;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_D_XOR;
  wire [0:0] CLBLM_R_X103Y124_SLICE_X163Y124_SR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A5Q;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_AMUX;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_AO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_AQ;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_A_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_BO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_BQ;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_B_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C5Q;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CLK;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CMUX;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_CQ;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_C_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_DO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_DO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_D_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X162Y125_SR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_AO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_AO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_AQ;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_A_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B5Q;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_BMUX;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_BO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_BO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_BQ;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_B_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C5Q;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CLK;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CMUX;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_CQ;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_C_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D1;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D2;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D3;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D4;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_DO5;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_DO6;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D_CY;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_D_XOR;
  wire [0:0] CLBLM_R_X103Y125_SLICE_X163Y125_SR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_AO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_AO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_AQ;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_A_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B5Q;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_BMUX;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_BO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_BO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_BQ;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_B_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_CLK;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_CO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_CO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_C_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_DO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_DO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_D_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X162Y126_SR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A5Q;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_AMUX;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_AO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_AO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_AQ;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_A_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_BO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_BO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_B_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_CLK;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_CO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_CO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_C_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D1;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D2;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D3;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D4;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_DO5;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_DO6;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D_CY;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_D_XOR;
  wire [0:0] CLBLM_R_X103Y126_SLICE_X163Y126_SR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_AO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_AO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_AQ;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_A_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_BO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_BO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_B_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_CLK;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_CO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_CO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_C_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_DO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_DO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_D_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X162Y127_SR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_AO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_AO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_A_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_BO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_BO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_B_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_CO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_CO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_C_XOR;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D1;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D2;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D3;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D4;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_DO5;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_DO6;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D_CY;
  wire [0:0] CLBLM_R_X103Y127_SLICE_X163Y127_D_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_AO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_AO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_A_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_BO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_BO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_B_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_CO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_CO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_C_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_DO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_DO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X140Y114_D_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A5Q;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_AMUX;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_AO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_AO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_AQ;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_A_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B5Q;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_BMUX;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_BO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_BO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_BQ;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_B_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_CLK;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_CO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_CO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_C_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D1;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D2;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D3;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D4;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_DO5;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_DO6;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D_CY;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_D_XOR;
  wire [0:0] CLBLM_R_X89Y114_SLICE_X141Y114_SR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A5Q;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_AMUX;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_AO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_AO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_AQ;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_AX;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_A_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_BMUX;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_BO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_BO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_B_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C5Q;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_CLK;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_CMUX;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_CO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_CO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_CQ;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_C_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_DO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_DO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_D_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X140Y115_SR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A5Q;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_AMUX;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_AO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_AO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_AQ;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_A_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B5Q;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_BMUX;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_BO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_BO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_BQ;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_B_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_CLK;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_CO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_CO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_CQ;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_C_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D1;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D2;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D3;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D4;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_DO5;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_DO6;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D_CY;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_D_XOR;
  wire [0:0] CLBLM_R_X89Y115_SLICE_X141Y115_SR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A5Q;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_AMUX;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_AO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_AO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_AQ;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_A_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B5Q;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_BMUX;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_BO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_BO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_BQ;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_BX;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_B_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_CLK;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_CO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_CO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_C_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_DO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_DO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_D_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X140Y116_SR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_AMUX;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_AO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_AO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_A_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B5Q;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_BMUX;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_BO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_BO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_BQ;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_B_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C5Q;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_CLK;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_CMUX;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_CO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_CO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_CQ;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_C_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D1;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D2;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D3;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D4;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_DO5;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_DO6;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D_CY;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_D_XOR;
  wire [0:0] CLBLM_R_X89Y116_SLICE_X141Y116_SR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A5Q;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_AMUX;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_AO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_AO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_AQ;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_A_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_BO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_BO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_BQ;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_B_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C5Q;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_CLK;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_CMUX;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_CO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_CO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_CQ;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_C_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_DO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_DO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_D_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X140Y117_SR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A5Q;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_AMUX;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_AO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_AO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_AQ;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_AX;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_A_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_BMUX;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_BO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_BO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_B_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C5Q;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_CLK;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_CMUX;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_CO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_CO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_CQ;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_C_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D1;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D2;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D3;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D4;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_DO5;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_DO6;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D_CY;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_D_XOR;
  wire [0:0] CLBLM_R_X89Y117_SLICE_X141Y117_SR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A5Q;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_AMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_AO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_AO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_AQ;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_A_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B5Q;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_BMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_BO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_BO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_BQ;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_BX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_B_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_CLK;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_CMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_CO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_CO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_C_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D5Q;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_DMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_DO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_DO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_DQ;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_D_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X140Y118_SR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A5Q;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_AMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_AO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_AO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_AQ;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_AX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_A_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_BMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_BO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_BO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_B_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_CLK;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_CO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_CO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_CQ;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_C_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D1;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D2;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D3;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D4;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D5Q;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_DMUX;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_DO5;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_DO6;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_DQ;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D_CY;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_D_XOR;
  wire [0:0] CLBLM_R_X89Y118_SLICE_X141Y118_SR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A5Q;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_AMUX;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_AO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_AO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_AQ;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_A_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B5Q;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_BMUX;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_BO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_BO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_BQ;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_B_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_CLK;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_CO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_CO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_C_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_DO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_DO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_D_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X140Y119_SR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A5Q;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_AMUX;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_AO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_AO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_AQ;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_AX;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_A_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_BMUX;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_BO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_BO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_B_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C5Q;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_CLK;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_CMUX;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_CO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_CO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_CQ;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_C_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D1;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D2;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D3;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D4;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_DO5;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_DO6;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D_CY;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_D_XOR;
  wire [0:0] CLBLM_R_X89Y119_SLICE_X141Y119_SR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A5Q;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_AMUX;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_AO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_AO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_AQ;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_AX;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_A_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_BMUX;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_BO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_BO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_B_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_CLK;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_CO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_CO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_CQ;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_C_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_DO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_DO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_D_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X140Y120_SR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A5Q;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_AMUX;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_AO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_AO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_AQ;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_A_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_BO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_BO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_BQ;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_B_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C5Q;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_CLK;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_CMUX;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_CO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_CO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_CQ;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_C_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D1;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D2;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D3;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D4;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_DO5;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_DO6;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D_CY;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_D_XOR;
  wire [0:0] CLBLM_R_X89Y120_SLICE_X141Y120_SR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A5Q;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_AMUX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_AO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_AO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_AQ;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_AX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_A_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_BMUX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_BO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_BO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_B_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C5Q;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_CLK;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_CMUX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_CO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_CO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_CQ;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_C_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_DO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_DO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_D_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X140Y121_SR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A5Q;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_AMUX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_AO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_AO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_AQ;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_AX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_A_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_BMUX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_BO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_BO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_B_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C5Q;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_CLK;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_CMUX;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_CO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_CO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_CQ;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_C_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D1;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D2;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D3;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D4;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_DO5;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_DO6;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D_CY;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_D_XOR;
  wire [0:0] CLBLM_R_X89Y121_SLICE_X141Y121_SR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A5Q;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_AMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_AO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_AO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_AQ;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_AX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_A_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_BMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_BO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_BO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_B_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C5Q;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_CLK;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_CMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_CO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_CO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_CQ;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_C_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_DO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_DO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_D_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X140Y122_SR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A5Q;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_AMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_AO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_AO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_AQ;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_A_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B5Q;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_BMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_BO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_BO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_BQ;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_BX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_B_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_CLK;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_CMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_CO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_CO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_C_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D1;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D2;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D3;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D4;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D5Q;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_DMUX;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_DO5;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_DO6;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_DQ;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D_CY;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_D_XOR;
  wire [0:0] CLBLM_R_X89Y122_SLICE_X141Y122_SR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A5Q;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_AMUX;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_AO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_AO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_AQ;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_AX;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_A_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_BMUX;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_BO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_BO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_B_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C5Q;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_CLK;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_CMUX;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_CO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_CO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_CQ;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_C_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_DO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_DO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_D_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X140Y123_SR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A5Q;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_AMUX;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_AO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_AO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_AQ;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_A_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_BO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_BO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_B_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_CLK;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_CO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_CO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_C_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D1;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D2;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D3;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D4;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_DO5;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_DO6;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D_CY;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_D_XOR;
  wire [0:0] CLBLM_R_X89Y123_SLICE_X141Y123_SR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A5Q;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_AMUX;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_AO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_AO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_AQ;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_A_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_BO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_BO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_BQ;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_B_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_CLK;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_CO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_CO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_CQ;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_C_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_DO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_DO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_D_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X140Y124_SR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A5Q;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_AMUX;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_AO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_AO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_AQ;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_A_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_BO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_BO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_BQ;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_B_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_CLK;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_CO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_CO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_C_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D1;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D2;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D3;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D4;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_DO5;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_DO6;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D_CY;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_D_XOR;
  wire [0:0] CLBLM_R_X89Y124_SLICE_X141Y124_SR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A5Q;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_AMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_AO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_AO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_AQ;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_A_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B5Q;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_BMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_BO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_BO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_BQ;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_BX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_B_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_CLK;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_CMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_CO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_CO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_C_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D5Q;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_DMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_DO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_DO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_DQ;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_D_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X140Y125_SR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A5Q;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_AMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_AO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_AO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_AQ;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_AX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_A_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_BMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_BO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_BO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_B_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C5Q;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_CLK;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_CMUX;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_CO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_CO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_CQ;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_C_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D1;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D2;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D3;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D4;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_DO5;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_DO6;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D_CY;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_D_XOR;
  wire [0:0] CLBLM_R_X89Y125_SLICE_X141Y125_SR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_AO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_AO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_AQ;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_A_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B5Q;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_BMUX;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_BO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_BO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_BQ;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_B_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_CLK;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_CO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_CO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_C_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_DO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_DO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_D_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X140Y126_SR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A5Q;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_AMUX;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_AO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_AO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_AQ;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_AX;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_A_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_BMUX;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_BO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_BO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_B_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C5Q;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_CLK;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_CMUX;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_CO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_CO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_CQ;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_C_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D1;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D2;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D3;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D4;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_DO5;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_DO6;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D_CY;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_D_XOR;
  wire [0:0] CLBLM_R_X89Y126_SLICE_X141Y126_SR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_AO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_AO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_A_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_BO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_BO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_B_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_CO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_CO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_C_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_DO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_DO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X140Y127_D_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A5Q;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_AMUX;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_AO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_AO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_AQ;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_A_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_BO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_BO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_B_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_CLK;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_CO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_CO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_C_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D1;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D2;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D3;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D4;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_DO5;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_DO6;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D_CY;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_D_XOR;
  wire [0:0] CLBLM_R_X89Y127_SLICE_X141Y127_SR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A5Q;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_AMUX;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_AO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_AO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_AQ;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_AX;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_A_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_BMUX;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_BO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_BO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_B_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C5Q;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_CLK;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_CMUX;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_CO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_CO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_CQ;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_C_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_DO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_DO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_D_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X140Y128_SR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A5Q;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_AMUX;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_AO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_AO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_AQ;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_A_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_BO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_BO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_B_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_CLK;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_CO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_CO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_C_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D1;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D2;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D3;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D4;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_DO5;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_DO6;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D_CY;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_D_XOR;
  wire [0:0] CLBLM_R_X89Y128_SLICE_X141Y128_SR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_AO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_AO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_AQ;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_A_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_BO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_BO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_B_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_CLK;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_CO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_CO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_C_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_DO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_DO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_D_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X140Y130_SR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A5Q;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_AMUX;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_AO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_AO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_AQ;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_A_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_BO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_BO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_BQ;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_B_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_CLK;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_CO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_CO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_C_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D1;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D2;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D3;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D4;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_DO5;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_DO6;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D_CY;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_D_XOR;
  wire [0:0] CLBLM_R_X89Y130_SLICE_X141Y130_SR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A5Q;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_AMUX;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_AO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_AO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_AQ;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_A_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_BO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_BO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_B_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_CLK;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_CO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_CO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_C_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_DO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_DO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_D_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X140Y131_SR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_AO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_AO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_A_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_BO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_BO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_B_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_CO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_CO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_C_XOR;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D1;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D2;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D3;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D4;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_DO5;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_DO6;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D_CY;
  wire [0:0] CLBLM_R_X89Y131_SLICE_X141Y131_D_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_AO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_AO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_A_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_BO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_BO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_B_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_CO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_CO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_C_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_DO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_DO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X146Y111_D_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A5Q;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_AMUX;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_AO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_AO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_AQ;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_A_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B5Q;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_BMUX;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_BO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_BO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_BQ;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_B_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_CLK;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_CO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_CO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_C_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D1;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D2;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D3;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D4;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_DO5;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_DO6;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D_CY;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_D_XOR;
  wire [0:0] CLBLM_R_X93Y111_SLICE_X147Y111_SR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A5Q;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_AMUX;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_AO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_AO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_AQ;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_A_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B5Q;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_BMUX;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_BO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_BO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_BQ;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_B_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_CLK;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_CO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_CO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_C_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_DO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_DO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_D_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X146Y112_SR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A5Q;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_AMUX;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_AO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_AO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_AQ;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_A_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B5Q;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_BMUX;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_BO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_BO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_BQ;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_B_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C5Q;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_CLK;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_CMUX;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_CO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_CO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_CQ;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_C_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D1;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D2;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D3;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D4;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_DO5;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_DO6;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D_CY;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_D_XOR;
  wire [0:0] CLBLM_R_X93Y112_SLICE_X147Y112_SR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A5Q;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_AMUX;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_AO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_AO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_AQ;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_A_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B5Q;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_BMUX;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_BO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_BO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_BQ;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_B_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_CLK;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_CO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_CO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_C_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_DO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_DO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_D_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X146Y113_SR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A5Q;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_AMUX;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_AO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_AO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_AQ;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_A_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B5Q;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_BMUX;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_BO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_BO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_BQ;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_B_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_CLK;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_CO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_CO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_C_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D1;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D2;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D3;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D4;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_DO5;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_DO6;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D_CY;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_D_XOR;
  wire [0:0] CLBLM_R_X93Y113_SLICE_X147Y113_SR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A5Q;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_AMUX;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_AO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_AO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_AQ;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_A_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B5Q;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_BMUX;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_BO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_BO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_BQ;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_B_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_CLK;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_CO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_CO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_C_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_DMUX;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_DO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_DO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_D_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X146Y114_SR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A5Q;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_AMUX;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_AO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_AO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_AQ;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_A_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B5Q;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_BMUX;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_BO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_BO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_BQ;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_B_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_CLK;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_CO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_CO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_C_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D1;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D2;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D3;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D4;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_DO5;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_DO6;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D_CY;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_D_XOR;
  wire [0:0] CLBLM_R_X93Y114_SLICE_X147Y114_SR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A5Q;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_AMUX;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_AO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_AO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_AQ;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_A_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B5Q;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_BMUX;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_BO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_BO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_BQ;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_B_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_CLK;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_CO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_CO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_C_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_DO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_DO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_D_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X146Y115_SR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A5Q;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_AMUX;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_AO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_AO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_AQ;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_A_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B5Q;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_BMUX;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_BO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_BO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_BQ;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_B_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_CLK;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_CMUX;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_CO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_CO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_C_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D1;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D2;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D3;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D4;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_DO5;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_DO6;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D_CY;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_D_XOR;
  wire [0:0] CLBLM_R_X93Y115_SLICE_X147Y115_SR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A5Q;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_AMUX;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_AO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_AO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_AQ;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_A_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B5Q;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_BMUX;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_BO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_BO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_BQ;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_B_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_CLK;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_CO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_CO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_C_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_DO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_DO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_D_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X146Y116_SR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A5Q;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_AMUX;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_AO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_AO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_AQ;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_A_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B5Q;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_BMUX;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_BO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_BO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_BQ;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_B_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_CLK;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_CO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_CO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_C_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D1;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D2;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D3;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D4;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_DO5;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_DO6;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D_CY;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_D_XOR;
  wire [0:0] CLBLM_R_X93Y116_SLICE_X147Y116_SR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A5Q;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_AMUX;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_AO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_AO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_AQ;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_A_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B5Q;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_BMUX;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_BO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_BO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_BQ;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_B_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_CLK;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_CO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_CO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_C_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_DO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_DO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_D_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X146Y117_SR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_AO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_AO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_A_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_BO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_BO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_B_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_CO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_CO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_C_XOR;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D1;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D2;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D3;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D4;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_DO5;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_DO6;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D_CY;
  wire [0:0] CLBLM_R_X93Y117_SLICE_X147Y117_D_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_AO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_AO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_A_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_BO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_BO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_B_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_CO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_CO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_C_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_DO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_DO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X146Y118_D_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A5Q;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_AMUX;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_AO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_AO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_AQ;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_A_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B5Q;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_BMUX;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_BO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_BO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_BQ;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_B_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_CLK;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_CO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_CO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_C_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D1;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D2;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D3;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D4;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_DO5;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_DO6;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D_CY;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_D_XOR;
  wire [0:0] CLBLM_R_X93Y118_SLICE_X147Y118_SR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A5Q;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_AMUX;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_AO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_AO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_AQ;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_A_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B5Q;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_BMUX;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_BO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_BO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_BQ;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_B_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C5Q;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_CLK;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_CMUX;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_CO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_CO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_CQ;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_C_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_DO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_DO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_D_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X146Y119_SR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A5Q;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_AMUX;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_AO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_AO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_AQ;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_A_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B5Q;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_BMUX;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_BO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_BO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_BQ;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_B_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_CLK;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_CO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_CO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_C_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D1;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D2;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D3;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D4;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_DO5;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_DO6;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D_CY;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_D_XOR;
  wire [0:0] CLBLM_R_X93Y119_SLICE_X147Y119_SR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A5Q;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_AMUX;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_AO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_AO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_AQ;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_A_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B5Q;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_BMUX;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_BO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_BO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_BQ;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_B_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_CLK;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_CO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_CO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_C_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_DO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_DO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_D_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X146Y120_SR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A5Q;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_AMUX;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_AO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_AO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_AQ;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_A_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B5Q;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_BMUX;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_BO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_BO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_BQ;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_B_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C5Q;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_CLK;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_CMUX;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_CO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_CO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_CQ;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_C_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D1;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D2;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D3;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D4;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_DO5;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_DO6;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D_CY;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_D_XOR;
  wire [0:0] CLBLM_R_X93Y120_SLICE_X147Y120_SR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A5Q;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_AMUX;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_AO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_AO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_AQ;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_A_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_BO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_BO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_BQ;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_B_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_CLK;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_CO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_CO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_CQ;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_C_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_DO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_DO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_D_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X146Y121_SR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_AMUX;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_AO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_AO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_AQ;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_A_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B5Q;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_BMUX;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_BO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_BO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_BQ;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_B_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C5Q;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_CLK;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_CMUX;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_CO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_CO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_CQ;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_C_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D1;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D2;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D3;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D4;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_DO5;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_DO6;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D_CY;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_D_XOR;
  wire [0:0] CLBLM_R_X93Y121_SLICE_X147Y121_SR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A5Q;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_AMUX;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_AO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_AO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_AQ;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_A_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_BO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_BO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_B_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_CLK;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_CO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_CO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_C_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_DO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_DO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_D_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X146Y122_SR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A5Q;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AMUX;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AQ;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_AX;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_A_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_BMUX;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_BO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_B_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C5Q;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CLK;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CMUX;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_CQ;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_C_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D1;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D2;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D3;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D4;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_DO5;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_DO6;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D_CY;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_D_XOR;
  wire [0:0] CLBLM_R_X93Y122_SLICE_X147Y122_SR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_AO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_AO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_AQ;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_A_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B5Q;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_BMUX;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_BO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_BO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_BQ;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_B_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_CLK;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_CO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_CO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_CQ;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_CX;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_C_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_DO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_DO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_D_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X146Y123_SR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_AMUX;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_AO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_AO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_A_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B5Q;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_BMUX;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_BO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_BO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_BQ;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_B_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C5Q;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_CLK;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_CMUX;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_CO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_CO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_CQ;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_C_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D1;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D2;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D3;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D4;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_DO5;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_DO6;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D_CY;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_D_XOR;
  wire [0:0] CLBLM_R_X93Y123_SLICE_X147Y123_SR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A5Q;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_AMUX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_AO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_AO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_AQ;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_AX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_A_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_BMUX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_BO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_BO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_B_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C5Q;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_CLK;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_CMUX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_CO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_CO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_CQ;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_C_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_DO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_DO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_D_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X146Y124_SR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A5Q;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_AMUX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_AO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_AO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_AQ;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_A_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B5Q;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_BMUX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_BO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_BO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_BQ;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_B_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C5Q;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_CLK;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_CMUX;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_CO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_CO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_CQ;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_C_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D1;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D2;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D3;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D4;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_DO5;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_DO6;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D_CY;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_D_XOR;
  wire [0:0] CLBLM_R_X93Y124_SLICE_X147Y124_SR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A5Q;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_AMUX;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_AO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_AO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_AQ;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_AX;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_A_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_BMUX;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_BO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_BO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_B_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C5Q;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_CLK;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_CMUX;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_CO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_CO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_CQ;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_C_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_DO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_DO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_D_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X146Y125_SR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A5Q;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_AMUX;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_AO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_AO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_AQ;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_A_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_BO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_BO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_B_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_CLK;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_CO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_CO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_C_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D1;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D2;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D3;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D4;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_DO5;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_DO6;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D_CY;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_D_XOR;
  wire [0:0] CLBLM_R_X93Y125_SLICE_X147Y125_SR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A5Q;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_AMUX;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_AO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_AO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_AQ;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_A_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_BO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_BO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_BQ;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_B_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C5Q;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_CLK;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_CMUX;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_CO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_CO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_CQ;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_C_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_DO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_DO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_D_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X146Y126_SR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A5Q;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_AMUX;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_AO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_AO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_AQ;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_AX;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_A_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_BMUX;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_BO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_BO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_B_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C5Q;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_CLK;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_CMUX;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_CO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_CO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_CQ;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_C_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D1;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D2;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D3;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D4;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_DO5;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_DO6;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D_CY;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_D_XOR;
  wire [0:0] CLBLM_R_X93Y126_SLICE_X147Y126_SR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A5Q;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_AMUX;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_AO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_AO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_AQ;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_A_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_BO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_BO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_BQ;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_B_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_CLK;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_CO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_CO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_CQ;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_C_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_DO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_DO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_D_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X146Y127_SR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_AO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_AO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_A_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_BO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_BO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_B_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_CO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_CO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_C_XOR;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D1;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D2;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D3;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D4;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_DO5;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_DO6;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D_CY;
  wire [0:0] CLBLM_R_X93Y127_SLICE_X147Y127_D_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A5Q;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_AMUX;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_AO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_AO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_AQ;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_AX;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_A_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_BMUX;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_BO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_BO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_B_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C5Q;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_CLK;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_CMUX;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_CO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_CO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_CQ;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_C_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_DO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_DO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_D_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X146Y128_SR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A5Q;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_AMUX;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_AO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_AO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_AQ;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_A_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B5Q;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_BMUX;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_BO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_BO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_BQ;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_B_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_CLK;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_CO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_CO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_CQ;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_C_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D1;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D2;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D3;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D4;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_DO5;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_DO6;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_DQ;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D_CY;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_D_XOR;
  wire [0:0] CLBLM_R_X93Y128_SLICE_X147Y128_SR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A5Q;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_AMUX;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_AO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_AO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_AQ;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_A_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B5Q;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_BMUX;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_BO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_BO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_BQ;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_B_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_CLK;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_CO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_CO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_CQ;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_C_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_DO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_DO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_D_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X146Y129_SR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A5Q;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_AMUX;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_AO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_AO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_AQ;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_A_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_BO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_BO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_B_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_CLK;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_CO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_CO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_C_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D1;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D2;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D3;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D4;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_DO5;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_DO6;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D_CY;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_D_XOR;
  wire [0:0] CLBLM_R_X93Y129_SLICE_X147Y129_SR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A5Q;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_AMUX;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_AO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_AO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_AQ;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_A_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B5Q;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_BMUX;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_BO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_BO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_BQ;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_B_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_CLK;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_CO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_CO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_C_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_DO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_DO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_D_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X146Y130_SR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A5Q;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_AMUX;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_AO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_AO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_AQ;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_AX;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_A_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_BMUX;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_BO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_BO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_B_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C5Q;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_CLK;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_CMUX;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_CO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_CO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_CQ;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_C_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D1;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D2;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D3;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D4;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_DO5;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_DO6;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D_CY;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_D_XOR;
  wire [0:0] CLBLM_R_X93Y130_SLICE_X147Y130_SR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A5Q;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_AMUX;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_AO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_AO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_AQ;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_AX;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_A_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_BMUX;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_BO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_BO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_B_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C5Q;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_CLK;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_CMUX;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_CO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_CO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_CQ;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_C_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_DO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_DO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_D_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X146Y131_SR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A5Q;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_AMUX;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_AO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_AO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_AQ;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_A_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B5Q;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_BMUX;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_BO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_BO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_BQ;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_B_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_CLK;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_CO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_CO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_C_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D1;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D2;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D3;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D4;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_DO5;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_DO6;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D_CY;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_D_XOR;
  wire [0:0] CLBLM_R_X93Y131_SLICE_X147Y131_SR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A5Q;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_AMUX;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_AO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_AO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_AQ;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_A_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_BO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_BO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_B_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_CLK;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_CO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_CO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_C_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_DO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_DO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_D_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X146Y132_SR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_AO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_AO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_A_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_BO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_BO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_B_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_CO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_CO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_C_XOR;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D1;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D2;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D3;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D4;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_DO5;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_DO6;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D_CY;
  wire [0:0] CLBLM_R_X93Y132_SLICE_X147Y132_D_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A5Q;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_AMUX;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_AO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_AO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_AQ;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_AX;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_A_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_BMUX;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_BO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_BO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_B_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C5Q;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_CLK;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_CMUX;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_CO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_CO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_CQ;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_C_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_DO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_DO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_D_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X146Y133_SR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_AO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_AO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_A_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_BO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_BO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_B_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_CO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_CO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_C_XOR;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D1;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D2;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D3;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D4;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_DO5;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_DO6;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D_CY;
  wire [0:0] CLBLM_R_X93Y133_SLICE_X147Y133_D_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A5Q;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_AMUX;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_AO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_AO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_AQ;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_A_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B5Q;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_BMUX;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_BO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_BO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_BQ;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_B_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C5Q;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_CLK;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_CMUX;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_CO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_CO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_CQ;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_C_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_DO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_DO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_D_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X150Y111_SR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A5Q;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_AMUX;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_AO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_AO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_AQ;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_A_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B5Q;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_BMUX;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_BO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_BO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_BQ;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_B_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_CLK;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_CO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_CO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_C_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D1;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D2;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D3;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D4;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_DO5;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_DO6;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D_CY;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_D_XOR;
  wire [0:0] CLBLM_R_X95Y111_SLICE_X151Y111_SR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A5Q;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_AMUX;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_AO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_AO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_AQ;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_A_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B5Q;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_BMUX;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_BO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_BO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_BQ;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_B_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_CLK;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_CMUX;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_CO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_CO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_C_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_DO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_DO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_D_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X150Y112_SR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_AMUX;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_AO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_AO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_A_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_BO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_BO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_B_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_CO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_CO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_C_XOR;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D1;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D2;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D3;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D4;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_DO5;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_DO6;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D_CY;
  wire [0:0] CLBLM_R_X95Y112_SLICE_X151Y112_D_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A5Q;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_AMUX;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_AO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_AO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_AQ;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_A_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B5Q;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_BMUX;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_BO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_BO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_BQ;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_B_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_CLK;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_CO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_CO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_C_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_DO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_DO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_D_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X150Y113_SR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A5Q;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_AMUX;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_AO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_AO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_AQ;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_A_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B5Q;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_BMUX;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_BO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_BO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_BQ;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_B_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_CLK;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_CO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_CO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_C_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D1;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D2;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D3;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D4;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_DO5;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_DO6;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D_CY;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_D_XOR;
  wire [0:0] CLBLM_R_X95Y113_SLICE_X151Y113_SR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A5Q;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_AMUX;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_AO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_AO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_AQ;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_A_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B5Q;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_BMUX;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_BO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_BO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_BQ;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_B_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C5Q;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_CLK;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_CMUX;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_CO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_CO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_CQ;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_C_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_DO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_DO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_D_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X150Y114_SR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_AO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_AO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_A_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_BO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_BO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_B_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_CO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_CO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_C_XOR;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D1;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D2;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D3;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D4;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_DO5;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_DO6;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D_CY;
  wire [0:0] CLBLM_R_X95Y114_SLICE_X151Y114_D_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A5Q;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_AMUX;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_AO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_AO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_AQ;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_A_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B5Q;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_BMUX;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_BO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_BO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_BQ;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_B_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C5Q;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_CLK;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_CMUX;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_CO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_CO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_CQ;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_C_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_DMUX;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_DO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_DO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_D_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X150Y115_SR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_AO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_AO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_A_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_BO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_BO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_B_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_CO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_CO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_C_XOR;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D1;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D2;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D3;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D4;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_DO5;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_DO6;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D_CY;
  wire [0:0] CLBLM_R_X95Y115_SLICE_X151Y115_D_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A5Q;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_AMUX;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_AO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_AO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_AQ;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_A_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_BO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_BO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_B_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_CLK;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_CO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_CO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_C_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_DO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_DO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_D_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X150Y116_SR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A5Q;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_AMUX;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_AO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_AO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_AQ;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_A_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_BO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_BO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_B_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_CLK;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_CO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_CO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_C_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D1;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D2;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D3;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D4;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_DO5;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_DO6;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D_CY;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_D_XOR;
  wire [0:0] CLBLM_R_X95Y116_SLICE_X151Y116_SR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A5Q;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_AMUX;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_AO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_AO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_AQ;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_A_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B5Q;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_BMUX;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_BO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_BO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_BQ;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_B_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C5Q;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_CLK;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_CMUX;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_CO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_CO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_CQ;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_C_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_DO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_DO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_D_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X150Y117_SR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_AO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_AO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_A_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_BO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_BO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_B_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_CO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_CO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_C_XOR;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D1;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D2;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D3;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D4;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_DO5;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_DO6;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D_CY;
  wire [0:0] CLBLM_R_X95Y117_SLICE_X151Y117_D_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A5Q;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_AMUX;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_AO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_AO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_AQ;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_A_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B5Q;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_BMUX;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_BO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_BO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_BQ;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_B_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C5Q;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_CLK;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_CMUX;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_CO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_CO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_CQ;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_C_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_DMUX;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_DO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_DO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_D_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X150Y118_SR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A5Q;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_AMUX;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_AO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_AO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_AQ;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_A_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B5Q;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_BMUX;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_BO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_BO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_BQ;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_B_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_CLK;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_CO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_CO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_C_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D1;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D2;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D3;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D4;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_DO5;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_DO6;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D_CY;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_D_XOR;
  wire [0:0] CLBLM_R_X95Y118_SLICE_X151Y118_SR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A5Q;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_AMUX;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_AO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_AO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_AQ;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_A_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B5Q;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_BMUX;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_BO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_BO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_BQ;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_B_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C5Q;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_CLK;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_CMUX;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_CO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_CO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_CQ;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_C_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_DO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_DO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_D_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X150Y119_SR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_AO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_AO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_A_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_BO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_BO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_B_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_CO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_CO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_C_XOR;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D1;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D2;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D3;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D4;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_DO5;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_DO6;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D_CY;
  wire [0:0] CLBLM_R_X95Y119_SLICE_X151Y119_D_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A5Q;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_AMUX;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_AO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_AO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_AQ;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_A_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B5Q;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_BMUX;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_BO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_BO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_BQ;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_B_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_CLK;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_CO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_CO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_C_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_DO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_DO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_D_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X150Y120_SR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A5Q;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_AMUX;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_AO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_AO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_AQ;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_A_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B5Q;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_BMUX;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_BO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_BO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_BQ;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_B_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_CLK;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_CO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_CO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_C_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D1;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D2;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D3;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D4;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_DO5;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_DO6;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D_CY;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_D_XOR;
  wire [0:0] CLBLM_R_X95Y120_SLICE_X151Y120_SR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A5Q;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_AMUX;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_AO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_AO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_AQ;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_A_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_BO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_BO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_B_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_CLK;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_CO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_CO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_C_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_DO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_DO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_D_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X150Y121_SR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A5Q;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_AMUX;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_AO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_AO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_AQ;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_A_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B5Q;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_BMUX;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_BO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_BO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_BQ;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_B_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_CLK;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_CMUX;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_CO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_CO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_C_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D1;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D2;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D3;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D4;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_DO5;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_DO6;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D_CY;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_D_XOR;
  wire [0:0] CLBLM_R_X95Y121_SLICE_X151Y121_SR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A5Q;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_AMUX;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_AO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_AO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_AQ;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_A_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B5Q;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_BMUX;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_BO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_BO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_BQ;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_B_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C5Q;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_CLK;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_CMUX;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_CO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_CO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_CQ;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_C_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_DO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_DO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_D_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X150Y122_SR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_AO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_AO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_A_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_BO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_BO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_B_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_CO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_CO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_C_XOR;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D1;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D2;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D3;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D4;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_DO5;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_DO6;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D_CY;
  wire [0:0] CLBLM_R_X95Y122_SLICE_X151Y122_D_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A5Q;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_AMUX;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_AO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_AO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_AQ;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_A_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B5Q;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_BMUX;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_BO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_BO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_BQ;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_B_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_CLK;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_CO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_CO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_C_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_DO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_DO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_D_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X150Y123_SR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A5Q;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_AMUX;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_AO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_AO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_AQ;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_A_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B5Q;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_BMUX;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_BO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_BO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_BQ;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_B_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_CLK;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_CO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_CO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_C_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D1;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D2;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D3;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D4;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_DO5;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_DO6;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D_CY;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_D_XOR;
  wire [0:0] CLBLM_R_X95Y123_SLICE_X151Y123_SR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A5Q;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_AMUX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_AO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_AO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_AQ;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_A_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B5Q;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_BMUX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_BO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_BO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_BQ;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_B_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C5Q;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_CLK;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_CMUX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_CO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_CO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_CQ;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_C_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_DO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_DO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_D_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X150Y124_SR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A5Q;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_AMUX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_AO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_AO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_AQ;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_AX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_A_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_BMUX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_BO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_BO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_B_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C5Q;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_CLK;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_CMUX;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_CO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_CO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_CQ;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_C_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D1;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D2;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D3;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D4;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_DO5;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_DO6;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D_CY;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_D_XOR;
  wire [0:0] CLBLM_R_X95Y124_SLICE_X151Y124_SR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A5Q;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_AMUX;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_AO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_AO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_AQ;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_A_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B5Q;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_BMUX;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_BO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_BO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_BQ;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_BX;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_B_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_CLK;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_CMUX;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_CO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_CO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_C_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_DO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_DO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_D_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X150Y125_SR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A5Q;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_AMUX;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_AO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_AO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_AQ;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_A_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_BO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_BO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_B_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_CLK;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_CO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_CO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_C_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D1;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D2;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D3;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D4;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_DO5;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_DO6;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D_CY;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_D_XOR;
  wire [0:0] CLBLM_R_X95Y125_SLICE_X151Y125_SR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A5Q;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_AMUX;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_AO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_AO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_AQ;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_A_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B5Q;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_BMUX;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_BO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_BO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_BQ;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_B_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_CLK;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_CO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_CO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_C_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_DO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_DO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_D_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X150Y126_SR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A5Q;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_AMUX;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_AO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_AO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_AQ;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_A_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_BO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_BO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_B_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_CLK;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_CO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_CO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_C_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D1;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D2;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D3;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D4;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_DO5;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_DO6;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D_CY;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_D_XOR;
  wire [0:0] CLBLM_R_X95Y126_SLICE_X151Y126_SR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_AO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_AO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_AQ;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_A_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B5Q;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_BMUX;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_BO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_BO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_BQ;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_B_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_CLK;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_CO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_CO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_C_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_DO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_DO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_D_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X150Y128_SR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_AO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_AO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_A_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_BO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_BO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_B_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_CO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_CO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_C_XOR;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D1;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D2;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D3;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D4;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_DO5;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_DO6;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D_CY;
  wire [0:0] CLBLM_R_X95Y128_SLICE_X151Y128_D_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A5Q;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_AMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_AO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_AO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_AQ;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_AX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_A_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_BMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_BO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_BO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_B_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C5Q;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_CLK;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_CMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_CO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_CO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_CQ;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_C_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_DO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_DO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_D_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X150Y129_SR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A5Q;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_AMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_AO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_AO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_AQ;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_A_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B5Q;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_BMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_BO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_BO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_BQ;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_BX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_B_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_CLK;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_CMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_CO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_CO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_C_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D1;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D2;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D3;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D4;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D5Q;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_DMUX;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_DO5;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_DO6;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_DQ;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D_CY;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_D_XOR;
  wire [0:0] CLBLM_R_X95Y129_SLICE_X151Y129_SR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A5Q;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_AMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_AO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_AO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_AQ;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_AX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_A_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_BMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_BO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_BO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_B_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C5Q;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_CLK;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_CMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_CO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_CO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_CQ;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_C_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_DMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_DO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_DO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_D_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X150Y130_SR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A5Q;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_AMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_AO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_AO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_AQ;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_AX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_A_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_BMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_BO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_BO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_B_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C5Q;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_CLK;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_CMUX;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_CO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_CO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_CQ;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_C_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D1;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D2;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D3;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D4;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_DO5;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_DO6;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D_CY;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_D_XOR;
  wire [0:0] CLBLM_R_X95Y130_SLICE_X151Y130_SR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A5Q;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_AMUX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_AO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_AO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_AQ;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_A_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B5Q;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_BMUX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_BO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_BO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_BQ;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_B_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_CLK;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_CO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_CO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_CQ;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_C_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_DO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_DO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_D_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X150Y131_SR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A5Q;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_AMUX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_AO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_AO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_AQ;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_AX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_A_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_BMUX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_BO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_BO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_B_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C5Q;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_CLK;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_CMUX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_CO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_CO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_CQ;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_C_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D1;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D2;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D3;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D4;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D5Q;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_DMUX;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_DO5;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_DO6;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_DQ;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D_CY;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_D_XOR;
  wire [0:0] CLBLM_R_X95Y131_SLICE_X151Y131_SR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_AO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_AO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_AQ;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_A_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B5Q;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_BMUX;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_BO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_BO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_BQ;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_B_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C5Q;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_CLK;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_CMUX;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_CO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_CO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_CQ;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_C_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_DO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_DO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_D_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X150Y132_SR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A5Q;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_AMUX;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_AO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_AO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_AQ;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_A_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B5Q;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_BMUX;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_BO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_BO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_BQ;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_BX;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_B_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_CLK;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_CO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_CO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_CQ;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_C_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D1;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D2;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D3;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D4;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_DMUX;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_DO5;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_DO6;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D_CY;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_D_XOR;
  wire [0:0] CLBLM_R_X95Y132_SLICE_X151Y132_SR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A5Q;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_AMUX;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_AO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_AO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_AQ;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_A_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B5Q;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_BMUX;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_BO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_BO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_BQ;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_B_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_CLK;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_CMUX;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_CO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_CO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_C_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_DO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_DO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_D_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X152Y111_SR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A5Q;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_AMUX;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_AO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_AO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_AQ;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_A_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_BO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_BO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_B_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_CLK;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_CO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_CO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_C_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D1;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D2;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D3;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D4;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_DO5;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_DO6;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D_CY;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_D_XOR;
  wire [0:0] CLBLM_R_X97Y111_SLICE_X153Y111_SR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A5Q;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_AMUX;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_AO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_AO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_AQ;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_A_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B5Q;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_BMUX;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_BO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_BO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_BQ;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_B_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C5Q;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_CLK;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_CMUX;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_CO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_CO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_CQ;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_C_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_DO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_DO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_D_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X152Y112_SR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A5Q;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_AMUX;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_AO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_AO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_AQ;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_A_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B5Q;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_BMUX;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_BO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_BO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_BQ;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_B_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_CLK;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_CMUX;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_CO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_CO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_C_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D1;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D2;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D3;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D4;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_DO5;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_DO6;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D_CY;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_D_XOR;
  wire [0:0] CLBLM_R_X97Y112_SLICE_X153Y112_SR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A5Q;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_AMUX;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_AO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_AO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_AQ;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_A_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_BO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_BO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_B_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_CLK;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_CO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_CO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_C_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_DO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_DO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_D_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X152Y113_SR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_AO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_AO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_A_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_BO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_BO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_B_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_CO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_CO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_C_XOR;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D1;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D2;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D3;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D4;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_DO5;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_DO6;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D_CY;
  wire [0:0] CLBLM_R_X97Y113_SLICE_X153Y113_D_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A5Q;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_AMUX;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_AO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_AO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_AQ;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_A_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_BO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_BO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_B_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_CLK;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_CO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_CO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_C_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_DO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_DO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_D_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X152Y115_SR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A5Q;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_AMUX;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_AO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_AO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_AQ;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_A_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B5Q;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_BMUX;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_BO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_BO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_BQ;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_B_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_CLK;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_CO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_CO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_C_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D1;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D2;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D3;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D4;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_DO5;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_DO6;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D_CY;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_D_XOR;
  wire [0:0] CLBLM_R_X97Y115_SLICE_X153Y115_SR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A5Q;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_AMUX;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_AO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_AO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_AQ;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_A_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B5Q;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_BMUX;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_BO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_BO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_BQ;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_B_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_CLK;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_CMUX;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_CO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_CO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_C_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_DO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_DO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_D_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X152Y116_SR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A5Q;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_AMUX;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_AO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_AO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_AQ;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_A_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B5Q;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_BMUX;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_BO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_BO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_BQ;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_B_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C5Q;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_CLK;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_CMUX;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_CO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_CO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_CQ;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_C_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D1;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D2;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D3;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D4;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_DO5;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_DO6;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D_CY;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_D_XOR;
  wire [0:0] CLBLM_R_X97Y116_SLICE_X153Y116_SR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A5Q;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_AMUX;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_AO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_AO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_AQ;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_A_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B5Q;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_BMUX;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_BO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_BO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_BQ;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_BX;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_B_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_CLK;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_CO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_CO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_C_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_DO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_DO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_D_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X152Y117_SR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A5Q;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_AMUX;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_AO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_AO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_AQ;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_A_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_BO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_BO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_BQ;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_B_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C5Q;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_CLK;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_CMUX;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_CO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_CO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_CQ;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_C_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D1;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D2;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D3;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D4;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_DMUX;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_DO5;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_DO6;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D_CY;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_D_XOR;
  wire [0:0] CLBLM_R_X97Y117_SLICE_X153Y117_SR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A5Q;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_AMUX;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_AO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_AO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_AQ;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_AX;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_A_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_BMUX;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_BO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_BO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_B_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C5Q;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_CLK;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_CMUX;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_CO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_CO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_CQ;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_C_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_DO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_DO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_D_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X152Y118_SR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_AO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_AO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_AQ;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_A_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B5Q;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_BMUX;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_BO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_BO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_BQ;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_B_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C5Q;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_CLK;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_CMUX;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_CO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_CO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_CQ;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_C_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D1;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D2;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D3;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D4;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_DO5;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_DO6;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D_CY;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_D_XOR;
  wire [0:0] CLBLM_R_X97Y118_SLICE_X153Y118_SR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A5Q;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_AMUX;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_AO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_AO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_AQ;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_A_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B5Q;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_BMUX;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_BO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_BO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_BQ;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_B_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_CLK;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_CO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_CO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_CQ;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_C_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_DO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_DO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_D_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X152Y119_SR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A5Q;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_AMUX;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_AO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_AO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_AQ;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_A_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_BO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_BO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_BQ;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_B_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C5Q;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_CLK;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_CMUX;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_CO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_CO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_CQ;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_C_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D1;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D2;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D3;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D4;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_DO5;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_DO6;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D_CY;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_D_XOR;
  wire [0:0] CLBLM_R_X97Y119_SLICE_X153Y119_SR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A5Q;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_AMUX;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_AO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_AO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_AQ;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_A_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_BO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_BO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_BQ;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_B_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_CLK;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_CMUX;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_CO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_CO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_C_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_DO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_DO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_D_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X152Y120_SR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A5Q;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_AMUX;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_AO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_AO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_AQ;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_A_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B5Q;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_BMUX;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_BO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_BO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_BQ;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_B_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C5Q;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_CLK;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_CMUX;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_CO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_CO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_CQ;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_C_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D1;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D2;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D3;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D4;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D5Q;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_DMUX;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_DO5;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_DO6;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_DQ;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D_CY;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_D_XOR;
  wire [0:0] CLBLM_R_X97Y120_SLICE_X153Y120_SR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A5Q;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_AMUX;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_AO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_AO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_AQ;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_A_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B5Q;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_BMUX;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_BO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_BO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_BQ;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_B_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C5Q;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_CLK;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_CMUX;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_CO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_CO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_CQ;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_C_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_DO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_DO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_D_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X152Y121_SR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A5Q;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_AMUX;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_AO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_AO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_AQ;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_A_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B5Q;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_BMUX;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_BO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_BO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_BQ;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_B_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C5Q;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_CLK;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_CMUX;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_CO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_CO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_CQ;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_C_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D1;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D2;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D3;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D4;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_DO5;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_DO6;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D_CY;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_D_XOR;
  wire [0:0] CLBLM_R_X97Y121_SLICE_X153Y121_SR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A5Q;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_AMUX;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_AO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_AO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_AQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_A_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_BO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_BO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_BQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_B_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_CLK;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_CO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_CO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_CQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_C_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D5Q;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_DMUX;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_DO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_DO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_DQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_D_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X152Y122_SR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_AO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_AO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_AQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_A_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B5Q;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_BMUX;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_BO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_BO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_BQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_B_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C5Q;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_CLK;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_CMUX;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_CO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_CO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_CQ;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_C_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D1;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D2;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D3;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D4;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_DO5;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_DO6;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D_CY;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_D_XOR;
  wire [0:0] CLBLM_R_X97Y122_SLICE_X153Y122_SR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A5Q;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_AMUX;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_AO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_AO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_AQ;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_A_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B5Q;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_BMUX;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_BO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_BO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_BQ;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_B_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C5Q;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_CLK;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_CMUX;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_CO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_CO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_CQ;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_C_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_DO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_DO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_D_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X152Y123_SR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A5Q;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_AMUX;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_AO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_AO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_AQ;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_A_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B5Q;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_BMUX;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_BO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_BO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_BQ;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_B_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C5Q;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_CLK;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_CMUX;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_CO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_CO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_CQ;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_C_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D1;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D2;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D3;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D4;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_DO5;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_DO6;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D_CY;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_D_XOR;
  wire [0:0] CLBLM_R_X97Y123_SLICE_X153Y123_SR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A5Q;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_AMUX;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_AO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_AO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_AQ;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_A_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B5Q;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_BMUX;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_BO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_BO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_BQ;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_B_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_CLK;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_CO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_CO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_C_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_DO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_DO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_D_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X152Y124_SR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_AO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_AO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_A_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_BO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_BO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_B_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_CO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_CO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_C_XOR;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D1;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D2;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D3;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D4;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_DO5;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_DO6;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D_CY;
  wire [0:0] CLBLM_R_X97Y124_SLICE_X153Y124_D_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A5Q;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_AMUX;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_AO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_AO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_AQ;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_A_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B5Q;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_BMUX;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_BO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_BO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_BQ;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_B_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_CLK;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_CO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_CO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_C_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_DO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_DO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_D_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X152Y125_SR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A5Q;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_AMUX;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_AO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_AO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_AQ;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_A_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B5Q;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_BMUX;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_BO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_BO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_BQ;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_B_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_CLK;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_CO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_CO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_C_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D1;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D2;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D3;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D4;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_DO5;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_DO6;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D_CY;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_D_XOR;
  wire [0:0] CLBLM_R_X97Y125_SLICE_X153Y125_SR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A5Q;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_AMUX;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_AO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_AO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_AQ;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_A_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B5Q;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_BMUX;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_BO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_BO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_BQ;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_B_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_CLK;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_CO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_CO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_C_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_DO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_DO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_D_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X152Y126_SR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_AO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_AO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_AQ;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_A_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B5Q;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_BMUX;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_BO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_BO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_BQ;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_B_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C5Q;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_CLK;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_CMUX;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_CO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_CO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_CQ;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_C_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D1;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D2;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D3;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D4;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_DO5;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_DO6;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D_CY;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_D_XOR;
  wire [0:0] CLBLM_R_X97Y126_SLICE_X153Y126_SR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A5Q;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_AMUX;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_AO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_AO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_AQ;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_A_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B5Q;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_BMUX;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_BO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_BO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_BQ;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_B_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_CLK;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_CMUX;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_CO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_CO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_C_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_DO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_DO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_D_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X152Y127_SR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A5Q;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_AMUX;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_AO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_AO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_AQ;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_A_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_BO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_BO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_BQ;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_B_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_CLK;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_CO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_CO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_C_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D1;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D2;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D3;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D4;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_DO5;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_DO6;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D_CY;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_D_XOR;
  wire [0:0] CLBLM_R_X97Y127_SLICE_X153Y127_SR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_AO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_AO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_AQ;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_A_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_BO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_BO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_B_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_CLK;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_CO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_CO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_C_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_DO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_DO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_D_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X152Y128_SR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A5Q;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_AMUX;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_AO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_AO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_AQ;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_AX;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_A_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_BMUX;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_BO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_BO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_B_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C5Q;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_CLK;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_CMUX;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_CO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_CO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_CQ;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_C_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D1;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D2;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D3;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D4;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_DO5;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_DO6;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D_CY;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_D_XOR;
  wire [0:0] CLBLM_R_X97Y128_SLICE_X153Y128_SR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A5Q;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_AMUX;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_AO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_AO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_AQ;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_A_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B5Q;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_BMUX;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_BO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_BO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_BQ;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_B_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_CLK;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_CO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_CO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_CQ;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_C_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_DO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_DO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_D_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X152Y129_SR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_AO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_AO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_A_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_BO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_BO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_B_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_CO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_CO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_C_XOR;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D1;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D2;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D3;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D4;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_DO5;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_DO6;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D_CY;
  wire [0:0] CLBLM_R_X97Y129_SLICE_X153Y129_D_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_AO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_AO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_AQ;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_A_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B5Q;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_BMUX;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_BO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_BO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_BQ;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_B_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_CLK;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_CO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_CO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_C_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_DO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_DO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_D_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X152Y130_SR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A5Q;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_AMUX;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_AO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_AO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_AQ;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_A_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_BO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_BO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_B_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_CLK;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_CO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_CO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_C_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D1;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D2;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D3;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D4;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_DO5;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_DO6;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D_CY;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_D_XOR;
  wire [0:0] CLBLM_R_X97Y130_SLICE_X153Y130_SR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_AO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_AO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_AQ;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_A_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B5Q;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_BMUX;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_BO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_BO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_BQ;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_B_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_CLK;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_CO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_CO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_C_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_DO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_DO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_D_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X152Y131_SR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_AO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_AO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_AQ;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_A_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B5Q;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_BMUX;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_BO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_BO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_BQ;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_B_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C5Q;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_CLK;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_CMUX;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_CO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_CO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_CQ;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_C_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D1;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D2;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D3;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D4;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_DO5;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_DO6;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D_CY;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_D_XOR;
  wire [0:0] CLBLM_R_X97Y131_SLICE_X153Y131_SR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A5Q;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_AMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_AO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_AO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_AQ;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_A_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B5Q;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_BMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_BO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_BO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_BQ;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_BX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_B_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_CLK;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_CMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_CO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_CO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_C_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D5Q;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_DMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_DO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_DO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_DQ;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_D_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X152Y132_SR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A5Q;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_AMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_AO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_AO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_AQ;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_A_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B5Q;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_BMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_BO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_BO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_BQ;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_B_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C5Q;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_CLK;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_CMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_CO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_CO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_CQ;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_C_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D1;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D2;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D3;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D4;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_DMUX;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_DO5;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_DO6;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D_CY;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_D_XOR;
  wire [0:0] CLBLM_R_X97Y132_SLICE_X153Y132_SR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A5Q;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_AMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_AO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_AO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_AQ;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_AX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_A_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_BMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_BO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_BO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_B_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C5Q;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_CLK;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_CMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_CO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_CO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_CQ;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_C_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_DO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_DO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_D_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X152Y133_SR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A5Q;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_AMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_AO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_AO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_AQ;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_AX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_A_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_BMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_BO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_BO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_B_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C5Q;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_CLK;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_CMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_CO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_CO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_CQ;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_C_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D1;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D2;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D3;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D4;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_DMUX;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_DO5;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_DO6;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D_CY;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_D_XOR;
  wire [0:0] CLBLM_R_X97Y133_SLICE_X153Y133_SR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_O;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_T;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_T;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_T;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_T;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_T;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_O;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_T;
  wire [0:0] LIOB33_SING_X0Y249_IOB_X0Y249_O;
  wire [0:0] LIOB33_SING_X0Y249_IOB_X0Y249_T;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_T;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_O;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_T;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_T;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_T;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_T;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_T;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_T;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_T;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_T;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_T;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_T;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_T;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_T;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_T;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_T;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_T;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_T;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_T;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_T;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_T;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_T;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_T;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_T;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_T;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_T;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_T;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_T;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_T;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_T;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_T;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_T;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_T;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_T;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_T;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_T;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_T;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_T;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_T;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_T;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_T;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_T;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_T;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_T;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_T;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_T;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_T;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_T;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_T;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_T;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_T;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_T;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_T;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_T;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_T;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_T;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_T;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_T;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_T;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_T;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_T;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_T;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_T;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_T;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_T;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_T;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_T;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_T;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_T;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_T;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_T;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_T;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_T;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_T;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_T;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_T;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_T;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_T;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_T;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_T;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_T;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_T;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_T;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_T;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_T;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_T;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_T;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_T;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_T;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_T;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_T;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_T;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_T;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_T;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_T;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_T;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_T;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_T;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_T;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_T;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y201_O;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y201_T;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y202_O;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y202_T;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y203_O;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y203_T;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y204_O;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y204_T;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y205_O;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y205_T;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y206_O;
  wire [0:0] LIOB33_X0Y205_IOB_X0Y206_T;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y207_O;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y207_T;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y208_O;
  wire [0:0] LIOB33_X0Y207_IOB_X0Y208_T;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y209_O;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y209_T;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y210_O;
  wire [0:0] LIOB33_X0Y209_IOB_X0Y210_T;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y211_O;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y211_T;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y212_O;
  wire [0:0] LIOB33_X0Y211_IOB_X0Y212_T;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y213_O;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y213_T;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y214_O;
  wire [0:0] LIOB33_X0Y213_IOB_X0Y214_T;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y215_O;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y215_T;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y216_O;
  wire [0:0] LIOB33_X0Y215_IOB_X0Y216_T;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y217_O;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y217_T;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y218_O;
  wire [0:0] LIOB33_X0Y217_IOB_X0Y218_T;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y219_O;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y219_T;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y220_O;
  wire [0:0] LIOB33_X0Y219_IOB_X0Y220_T;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y221_O;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y221_T;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y222_O;
  wire [0:0] LIOB33_X0Y221_IOB_X0Y222_T;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y223_O;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y223_T;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y224_O;
  wire [0:0] LIOB33_X0Y223_IOB_X0Y224_T;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y225_O;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y225_T;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y226_O;
  wire [0:0] LIOB33_X0Y225_IOB_X0Y226_T;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y227_O;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y227_T;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y228_O;
  wire [0:0] LIOB33_X0Y227_IOB_X0Y228_T;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y229_O;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y229_T;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y230_O;
  wire [0:0] LIOB33_X0Y229_IOB_X0Y230_T;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y231_O;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y231_T;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y232_O;
  wire [0:0] LIOB33_X0Y231_IOB_X0Y232_T;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y233_O;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y233_T;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y234_O;
  wire [0:0] LIOB33_X0Y233_IOB_X0Y234_T;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y235_O;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y235_T;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y236_O;
  wire [0:0] LIOB33_X0Y235_IOB_X0Y236_T;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y237_O;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y237_T;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y238_O;
  wire [0:0] LIOB33_X0Y237_IOB_X0Y238_T;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y239_O;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y239_T;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y240_O;
  wire [0:0] LIOB33_X0Y239_IOB_X0Y240_T;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y241_O;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y241_T;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y242_O;
  wire [0:0] LIOB33_X0Y241_IOB_X0Y242_T;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y243_O;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y243_T;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y244_O;
  wire [0:0] LIOB33_X0Y243_IOB_X0Y244_T;
  wire [0:0] LIOB33_X0Y245_IOB_X0Y245_O;
  wire [0:0] LIOB33_X0Y245_IOB_X0Y245_T;
  wire [0:0] LIOB33_X0Y245_IOB_X0Y246_O;
  wire [0:0] LIOB33_X0Y245_IOB_X0Y246_T;
  wire [0:0] LIOB33_X0Y247_IOB_X0Y247_O;
  wire [0:0] LIOB33_X0Y247_IOB_X0Y247_T;
  wire [0:0] LIOB33_X0Y247_IOB_X0Y248_O;
  wire [0:0] LIOB33_X0Y247_IOB_X0Y248_T;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_T;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_T;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_T;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_T;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_O;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_T;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_O;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_T;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_T;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_T;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_T;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_T;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_T;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_T;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_T;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_T;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_O;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_T;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_O;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_T;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_O;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_T;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_T;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_T;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_T;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_O;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_T;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_O;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_T;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_O;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_T;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_O;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_T;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_O;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_T;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_O;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_T;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_O;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_T;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_O;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_T;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_O;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_T;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_O;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_T;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_T;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_T;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_O;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_T;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_T;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_O;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_T;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_O;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_T;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_O;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_T;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_O;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_T;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_O;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_T;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_O;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_T;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_O;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_T;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_O;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_T;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_O;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_T;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_O;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_T;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_O;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_T;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_O;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_T;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_O;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_T;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_O;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_T;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_O;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_T;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_O;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_T;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_O;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_T;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_O;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_T;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_D1;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_OQ;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_T1;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_TQ;
  wire [0:0] LIOI3_SING_X0Y249_OLOGIC_X0Y249_D1;
  wire [0:0] LIOI3_SING_X0Y249_OLOGIC_X0Y249_OQ;
  wire [0:0] LIOI3_SING_X0Y249_OLOGIC_X0Y249_T1;
  wire [0:0] LIOI3_SING_X0Y249_OLOGIC_X0Y249_TQ;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_D1;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_OQ;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_T1;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_TQ;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_D1;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_OQ;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_T1;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y201_D1;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y201_OQ;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y201_T1;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y201_TQ;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y202_D1;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y202_OQ;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y202_T1;
  wire [0:0] LIOI3_X0Y201_OLOGIC_X0Y202_TQ;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y203_D1;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y203_OQ;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y203_T1;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y203_TQ;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y204_D1;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y204_OQ;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y204_T1;
  wire [0:0] LIOI3_X0Y203_OLOGIC_X0Y204_TQ;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y205_D1;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y205_OQ;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y205_T1;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y205_TQ;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y206_D1;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y206_OQ;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y206_T1;
  wire [0:0] LIOI3_X0Y205_OLOGIC_X0Y206_TQ;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y209_D1;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y209_OQ;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y209_T1;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y209_TQ;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y210_D1;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y210_OQ;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y210_T1;
  wire [0:0] LIOI3_X0Y209_OLOGIC_X0Y210_TQ;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y211_D1;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y211_OQ;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y211_T1;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y211_TQ;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y212_D1;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y212_OQ;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y212_T1;
  wire [0:0] LIOI3_X0Y211_OLOGIC_X0Y212_TQ;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y215_D1;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y215_OQ;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y215_T1;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y215_TQ;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y216_D1;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y216_OQ;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y216_T1;
  wire [0:0] LIOI3_X0Y215_OLOGIC_X0Y216_TQ;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y217_D1;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y217_OQ;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y217_T1;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y217_TQ;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y218_D1;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y218_OQ;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y218_T1;
  wire [0:0] LIOI3_X0Y217_OLOGIC_X0Y218_TQ;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y221_D1;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y221_OQ;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y221_T1;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y221_TQ;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y222_D1;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y222_OQ;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y222_T1;
  wire [0:0] LIOI3_X0Y221_OLOGIC_X0Y222_TQ;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y223_D1;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y223_OQ;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y223_T1;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y223_TQ;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y224_D1;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y224_OQ;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y224_T1;
  wire [0:0] LIOI3_X0Y223_OLOGIC_X0Y224_TQ;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y225_D1;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y225_OQ;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y225_T1;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y225_TQ;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y226_D1;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y226_OQ;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y226_T1;
  wire [0:0] LIOI3_X0Y225_OLOGIC_X0Y226_TQ;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y227_D1;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y227_OQ;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y227_T1;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y227_TQ;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y228_D1;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y228_OQ;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y228_T1;
  wire [0:0] LIOI3_X0Y227_OLOGIC_X0Y228_TQ;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y229_D1;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y229_OQ;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y229_T1;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y229_TQ;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y230_D1;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y230_OQ;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y230_T1;
  wire [0:0] LIOI3_X0Y229_OLOGIC_X0Y230_TQ;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y233_D1;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y233_OQ;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y233_T1;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y233_TQ;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y234_D1;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y234_OQ;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y234_T1;
  wire [0:0] LIOI3_X0Y233_OLOGIC_X0Y234_TQ;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y235_D1;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y235_OQ;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y235_T1;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y235_TQ;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y236_D1;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y236_OQ;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y236_T1;
  wire [0:0] LIOI3_X0Y235_OLOGIC_X0Y236_TQ;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y239_D1;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y239_OQ;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y239_T1;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y239_TQ;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y240_D1;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y240_OQ;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y240_T1;
  wire [0:0] LIOI3_X0Y239_OLOGIC_X0Y240_TQ;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y241_D1;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y241_OQ;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y241_T1;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y241_TQ;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y242_D1;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y242_OQ;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y242_T1;
  wire [0:0] LIOI3_X0Y241_OLOGIC_X0Y242_TQ;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y245_D1;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y245_OQ;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y245_T1;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y245_TQ;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y246_D1;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y246_OQ;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y246_T1;
  wire [0:0] LIOI3_X0Y245_OLOGIC_X0Y246_TQ;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y247_D1;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y247_OQ;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y247_T1;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y247_TQ;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y248_D1;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y248_OQ;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y248_T1;
  wire [0:0] LIOI3_X0Y247_OLOGIC_X0Y248_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_TQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_D1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_OQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_T1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_TQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_D1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_OQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_T1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_TQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_D1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_OQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_T1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_TQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_D1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_OQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_T1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_TQ;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y5_D1;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y5_OQ;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y5_T1;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y5_TQ;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y6_D1;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y6_OQ;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y6_T1;
  wire [0:0] LIOI3_X0Y5_OLOGIC_X0Y6_TQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_D1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_OQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_T1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_TQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_D1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_OQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_T1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_D1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_OQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_T1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y67_TQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_D1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_OQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_T1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_TQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_D1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_OQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_T1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y71_TQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_D1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_OQ;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_T1;
  wire [0:0] LIOI3_X0Y71_OLOGIC_X0Y72_TQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_D1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_OQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_T1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y73_TQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_D1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_OQ;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_T1;
  wire [0:0] LIOI3_X0Y73_OLOGIC_X0Y74_TQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_D1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_OQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_T1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y75_TQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_D1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_OQ;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_T1;
  wire [0:0] LIOI3_X0Y75_OLOGIC_X0Y76_TQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_D1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_OQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_T1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y77_TQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_D1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_OQ;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_T1;
  wire [0:0] LIOI3_X0Y77_OLOGIC_X0Y78_TQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y79_TQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_D1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_OQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_T1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y83_TQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_D1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_OQ;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_T1;
  wire [0:0] LIOI3_X0Y83_OLOGIC_X0Y84_TQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_D1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_OQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_T1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y85_TQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_D1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_OQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_T1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_TQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_D1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_OQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_T1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_TQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_D1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_OQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_T1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_TQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_D1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_OQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_T1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_TQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_D1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_OQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_T1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_TQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_D1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_OQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_T1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_TQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_D1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_OQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_T1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_TQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_D1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_OQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_T1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_TQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_D1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_OQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_T1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_T;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_T;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_T;
  wire [0:0] RIOB33_SING_X105Y99_IOB_X1Y99_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_T;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_T;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_T;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_T;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_T;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_T;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_T;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_T;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_T;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_T;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_T;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_T;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_T;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_T;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_T;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_T;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_T;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_T;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_T;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_T;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_T;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_T;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_T;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_T;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_T;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_T;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_T;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_T;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_T;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_T;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_T;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_T;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_T;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_T;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_T;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_T;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_T;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_T;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_T;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_T;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_T;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_T;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_T;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_T;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_T;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_T;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_T;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_T;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_T;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_T;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_T;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_T;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_T;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_T;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_T;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_T;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_T;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_T;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_T;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_T;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_T;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_T;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_T;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_T;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_T;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_T;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_T;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_T;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_T;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_T;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_T;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_T;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_T;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_T;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_T;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_T;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_T;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_I;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_T;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y92_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y93_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y94_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y95_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y96_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y97_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y98_O;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y78_D;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y78_O;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_TQ;


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X156Y111_AO5),
.Q(CLBLL_L_X100Y111_SLICE_X156Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X156Y111_BO5),
.Q(CLBLL_L_X100Y111_SLICE_X156Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X156Y111_AO6),
.Q(CLBLL_L_X100Y111_SLICE_X156Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X156Y111_BO6),
.Q(CLBLL_L_X100Y111_SLICE_X156Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_DLUT (
.I0(CLBLM_L_X98Y111_SLICE_X155Y111_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X100Y111_SLICE_X156Y111_BQ),
.I4(CLBLL_L_X100Y111_SLICE_X156Y111_B5Q),
.I5(CLBLM_R_X101Y111_SLICE_X158Y111_A5Q),
.O5(CLBLL_L_X100Y111_SLICE_X156Y111_DO5),
.O6(CLBLL_L_X100Y111_SLICE_X156Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1fbf15b51aba10b0)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y111_SLICE_X159Y111_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y111_SLICE_X156Y111_A5Q),
.I4(CLBLL_L_X100Y111_SLICE_X156Y111_DO6),
.I5(CLBLM_L_X98Y111_SLICE_X155Y111_DO6),
.O5(CLBLL_L_X100Y111_SLICE_X156Y111_CO5),
.O6(CLBLL_L_X100Y111_SLICE_X156Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y111_SLICE_X156Y111_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y111_SLICE_X155Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y111_SLICE_X156Y111_BO5),
.O6(CLBLL_L_X100Y111_SLICE_X156Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLL_L_X100Y111_SLICE_X156Y111_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y111_SLICE_X156Y111_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X100Y111_SLICE_X157Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y111_SLICE_X156Y111_AO5),
.O6(CLBLL_L_X100Y111_SLICE_X156Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X157Y111_AO5),
.Q(CLBLL_L_X100Y111_SLICE_X157Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X157Y111_BO5),
.Q(CLBLL_L_X100Y111_SLICE_X157Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X157Y111_CO5),
.Q(CLBLL_L_X100Y111_SLICE_X157Y111_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X157Y111_AO6),
.Q(CLBLL_L_X100Y111_SLICE_X157Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X157Y111_BO6),
.Q(CLBLL_L_X100Y111_SLICE_X157Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y111_SLICE_X157Y111_CO6),
.Q(CLBLL_L_X100Y111_SLICE_X157Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055e4e4aaffe4e4)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y111_SLICE_X152Y111_DO6),
.I2(CLBLM_R_X101Y111_SLICE_X158Y111_DO6),
.I3(CLBLM_R_X101Y111_SLICE_X159Y111_B5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X100Y111_SLICE_X157Y111_AQ),
.O5(CLBLL_L_X100Y111_SLICE_X157Y111_DO5),
.O6(CLBLL_L_X100Y111_SLICE_X157Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444cc0000cc)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_CLUT (
.I0(CLBLM_R_X101Y111_SLICE_X158Y111_CO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X100Y113_SLICE_X157Y113_A5Q),
.I4(CLBLM_L_X98Y111_SLICE_X154Y111_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y111_SLICE_X157Y111_CO5),
.O6(CLBLL_L_X100Y111_SLICE_X157Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc88884444)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_BLUT (
.I0(CLBLM_L_X98Y111_SLICE_X154Y111_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X100Y111_SLICE_X157Y111_DO6),
.I4(CLBLL_L_X100Y111_SLICE_X157Y111_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y111_SLICE_X157Y111_BO5),
.O6(CLBLL_L_X100Y111_SLICE_X157Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cc00cc00)
  ) CLBLL_L_X100Y111_SLICE_X157Y111_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X100Y115_SLICE_X156Y115_AQ),
.I4(CLBLL_L_X100Y111_SLICE_X157Y111_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y111_SLICE_X157Y111_AO5),
.O6(CLBLL_L_X100Y111_SLICE_X157Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y112_SLICE_X156Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y112_SLICE_X156Y112_AO5),
.Q(CLBLL_L_X100Y112_SLICE_X156Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y112_SLICE_X156Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y112_SLICE_X156Y112_AO6),
.Q(CLBLL_L_X100Y112_SLICE_X156Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y112_SLICE_X156Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y112_SLICE_X156Y112_DO5),
.O6(CLBLL_L_X100Y112_SLICE_X156Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLL_L_X100Y112_SLICE_X156Y112_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y112_SLICE_X156Y112_AQ),
.I2(1'b1),
.I3(CLBLL_L_X100Y112_SLICE_X156Y112_A5Q),
.I4(CLBLL_L_X100Y113_SLICE_X156Y113_A5Q),
.I5(CLBLM_L_X98Y112_SLICE_X154Y112_BQ),
.O5(CLBLL_L_X100Y112_SLICE_X156Y112_CO5),
.O6(CLBLL_L_X100Y112_SLICE_X156Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f77220a0a7722)
  ) CLBLL_L_X100Y112_SLICE_X156Y112_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y112_SLICE_X158Y112_B5Q),
.I2(CLBLL_L_X100Y111_SLICE_X156Y111_AQ),
.I3(CLBLM_R_X97Y112_SLICE_X152Y112_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X101Y112_SLICE_X158Y112_CO6),
.O5(CLBLL_L_X100Y112_SLICE_X156Y112_BO5),
.O6(CLBLL_L_X100Y112_SLICE_X156Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00c0c0c0c0)
  ) CLBLL_L_X100Y112_SLICE_X156Y112_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X100Y112_SLICE_X156Y112_AQ),
.I3(CLBLM_L_X98Y112_SLICE_X154Y112_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y112_SLICE_X156Y112_AO5),
.O6(CLBLL_L_X100Y112_SLICE_X156Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y112_SLICE_X157Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y112_SLICE_X157Y112_AO5),
.Q(CLBLL_L_X100Y112_SLICE_X157Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y112_SLICE_X157Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y112_SLICE_X157Y112_AO6),
.Q(CLBLL_L_X100Y112_SLICE_X157Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y112_SLICE_X157Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y112_SLICE_X157Y112_DO5),
.O6(CLBLL_L_X100Y112_SLICE_X157Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y112_SLICE_X157Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y112_SLICE_X157Y112_CO5),
.O6(CLBLL_L_X100Y112_SLICE_X157Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y112_SLICE_X157Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y112_SLICE_X157Y112_BO5),
.O6(CLBLL_L_X100Y112_SLICE_X157Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444cc0000cc)
  ) CLBLL_L_X100Y112_SLICE_X157Y112_ALUT (
.I0(CLBLL_L_X102Y112_SLICE_X160Y112_CO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X101Y112_SLICE_X158Y112_B5Q),
.I4(CLBLL_L_X100Y113_SLICE_X156Y113_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y112_SLICE_X157Y112_AO5),
.O6(CLBLL_L_X100Y112_SLICE_X157Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X156Y113_AO5),
.Q(CLBLL_L_X100Y113_SLICE_X156Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X156Y113_BO5),
.Q(CLBLL_L_X100Y113_SLICE_X156Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X156Y113_CO5),
.Q(CLBLL_L_X100Y113_SLICE_X156Y113_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X156Y113_AO6),
.Q(CLBLL_L_X100Y113_SLICE_X156Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X156Y113_BO6),
.Q(CLBLL_L_X100Y113_SLICE_X156Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X156Y113_CO6),
.Q(CLBLL_L_X100Y113_SLICE_X156Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_DLUT (
.I0(CLBLM_L_X98Y113_SLICE_X154Y113_AQ),
.I1(CLBLL_L_X100Y113_SLICE_X156Y113_AQ),
.I2(CLBLL_L_X100Y113_SLICE_X156Y113_BQ),
.I3(1'b1),
.I4(CLBLL_L_X100Y113_SLICE_X156Y113_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_DO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030f00000f0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y113_SLICE_X158Y113_CO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X100Y112_SLICE_X157Y112_A5Q),
.I4(CLBLL_L_X100Y113_SLICE_X156Y113_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_CO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y113_SLICE_X156Y113_BQ),
.I2(CLBLL_L_X100Y113_SLICE_X156Y113_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_BO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y112_SLICE_X156Y112_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X98Y113_SLICE_X154Y113_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_AO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X157Y113_AO5),
.Q(CLBLL_L_X100Y113_SLICE_X157Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y113_SLICE_X157Y113_AO6),
.Q(CLBLL_L_X100Y113_SLICE_X157Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_DO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_CO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5140d9c87362fbea)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X101Y112_SLICE_X159Y112_DO6),
.I3(CLBLM_L_X98Y110_SLICE_X154Y110_BO6),
.I4(CLBLL_L_X100Y115_SLICE_X156Y115_AQ),
.I5(CLBLL_L_X102Y113_SLICE_X161Y113_A5Q),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_BO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaa0a00a0a)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y114_SLICE_X154Y114_C5Q),
.I3(CLBLL_L_X100Y113_SLICE_X157Y113_BO6),
.I4(CLBLL_L_X100Y115_SLICE_X156Y115_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_AO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y114_SLICE_X156Y114_AO5),
.Q(CLBLL_L_X100Y114_SLICE_X156Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y114_SLICE_X156Y114_BO5),
.Q(CLBLL_L_X100Y114_SLICE_X156Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y114_SLICE_X156Y114_AO6),
.Q(CLBLL_L_X100Y114_SLICE_X156Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y114_SLICE_X156Y114_BO6),
.Q(CLBLL_L_X100Y114_SLICE_X156Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0afa0afa0c0cfcfc)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_DLUT (
.I0(CLBLM_R_X101Y113_SLICE_X159Y113_DO6),
.I1(CLBLM_L_X98Y114_SLICE_X154Y114_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y115_SLICE_X156Y115_A5Q),
.I4(CLBLL_L_X102Y114_SLICE_X160Y114_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y114_SLICE_X156Y114_DO5),
.O6(CLBLL_L_X100Y114_SLICE_X156Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f505f500c0cfcfc)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_CLUT (
.I0(CLBLL_L_X100Y114_SLICE_X156Y114_A5Q),
.I1(CLBLM_L_X94Y115_SLICE_X148Y115_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y115_SLICE_X155Y115_DO6),
.I4(CLBLL_L_X100Y114_SLICE_X156Y114_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y114_SLICE_X156Y114_CO5),
.O6(CLBLL_L_X100Y114_SLICE_X156Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y114_SLICE_X158Y114_CO6),
.I2(CLBLL_L_X100Y113_SLICE_X156Y113_C5Q),
.I3(CLBLM_L_X98Y115_SLICE_X155Y115_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y114_SLICE_X156Y114_BO5),
.O6(CLBLL_L_X100Y114_SLICE_X156Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X100Y114_SLICE_X156Y114_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y114_SLICE_X156Y114_A5Q),
.I2(CLBLM_L_X98Y112_SLICE_X154Y112_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y114_SLICE_X156Y114_AO5),
.O6(CLBLL_L_X100Y114_SLICE_X156Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y114_SLICE_X157Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y114_SLICE_X157Y114_DO5),
.O6(CLBLL_L_X100Y114_SLICE_X157Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y114_SLICE_X157Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y114_SLICE_X157Y114_CO5),
.O6(CLBLL_L_X100Y114_SLICE_X157Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y114_SLICE_X157Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y114_SLICE_X157Y114_BO5),
.O6(CLBLL_L_X100Y114_SLICE_X157Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y114_SLICE_X157Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y114_SLICE_X157Y114_AO5),
.O6(CLBLL_L_X100Y114_SLICE_X157Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X156Y115_AO5),
.Q(CLBLL_L_X100Y115_SLICE_X156Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X156Y115_BO5),
.Q(CLBLL_L_X100Y115_SLICE_X156Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X156Y115_CO5),
.Q(CLBLL_L_X100Y115_SLICE_X156Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X156Y115_AO6),
.Q(CLBLL_L_X100Y115_SLICE_X156Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X156Y115_BO6),
.Q(CLBLL_L_X100Y115_SLICE_X156Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X156Y115_CO6),
.Q(CLBLL_L_X100Y115_SLICE_X156Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff550033f033f0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_DLUT (
.I0(CLBLL_L_X100Y116_SLICE_X156Y116_AQ),
.I1(CLBLL_L_X102Y115_SLICE_X160Y115_A5Q),
.I2(CLBLM_L_X98Y115_SLICE_X154Y115_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y116_SLICE_X158Y116_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y115_SLICE_X156Y115_DO5),
.O6(CLBLL_L_X100Y115_SLICE_X156Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0c030c030)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y116_SLICE_X155Y116_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y115_SLICE_X153Y115_B5Q),
.I4(CLBLL_L_X100Y115_SLICE_X156Y115_DO6),
.I5(1'b1),
.O5(CLBLL_L_X100Y115_SLICE_X156Y115_CO5),
.O6(CLBLL_L_X100Y115_SLICE_X156Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222aa0000aa)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y114_SLICE_X156Y114_DO6),
.I2(1'b1),
.I3(CLBLM_L_X98Y114_SLICE_X154Y114_B5Q),
.I4(CLBLL_L_X100Y115_SLICE_X156Y115_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y115_SLICE_X156Y115_BO5),
.O6(CLBLL_L_X100Y115_SLICE_X156Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X100Y115_SLICE_X156Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y115_SLICE_X156Y115_A5Q),
.I2(CLBLL_L_X100Y116_SLICE_X156Y116_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y115_SLICE_X156Y115_AO5),
.O6(CLBLL_L_X100Y115_SLICE_X156Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X157Y115_BO5),
.Q(CLBLL_L_X100Y115_SLICE_X157Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X157Y115_AO6),
.Q(CLBLL_L_X100Y115_SLICE_X157Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y115_SLICE_X157Y115_BO6),
.Q(CLBLL_L_X100Y115_SLICE_X157Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699696696996)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_DLUT (
.I0(CLBLL_L_X100Y115_SLICE_X157Y115_BQ),
.I1(CLBLM_R_X101Y115_SLICE_X158Y115_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y115_SLICE_X157Y115_AQ),
.I4(CLBLL_L_X100Y115_SLICE_X157Y115_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y115_SLICE_X157Y115_DO5),
.O6(CLBLL_L_X100Y115_SLICE_X157Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969699696)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_CLUT (
.I0(CLBLL_L_X100Y115_SLICE_X157Y115_BQ),
.I1(CLBLL_L_X100Y115_SLICE_X157Y115_AQ),
.I2(CLBLM_R_X101Y115_SLICE_X158Y115_A5Q),
.I3(CLBLL_L_X102Y117_SLICE_X161Y117_A5Q),
.I4(CLBLL_L_X100Y115_SLICE_X157Y115_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X100Y115_SLICE_X157Y115_CO5),
.O6(CLBLL_L_X100Y115_SLICE_X157Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y115_SLICE_X157Y115_BQ),
.I2(CLBLL_L_X100Y115_SLICE_X157Y115_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y115_SLICE_X157Y115_BO5),
.O6(CLBLL_L_X100Y115_SLICE_X157Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a8a8202020a820)
  ) CLBLL_L_X100Y115_SLICE_X157Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y117_SLICE_X154Y117_AO6),
.I3(CLBLL_L_X100Y115_SLICE_X157Y115_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X102Y117_SLICE_X161Y117_A5Q),
.O5(CLBLL_L_X100Y115_SLICE_X157Y115_AO5),
.O6(CLBLL_L_X100Y115_SLICE_X157Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X156Y116_AO5),
.Q(CLBLL_L_X100Y116_SLICE_X156Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X156Y116_BO5),
.Q(CLBLL_L_X100Y116_SLICE_X156Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X156Y116_AO6),
.Q(CLBLL_L_X100Y116_SLICE_X156Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X156Y116_BO6),
.Q(CLBLL_L_X100Y116_SLICE_X156Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_DLUT (
.I0(CLBLM_L_X98Y116_SLICE_X155Y116_AQ),
.I1(CLBLM_R_X101Y116_SLICE_X158Y116_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X100Y116_SLICE_X156Y116_BQ),
.I4(CLBLL_L_X100Y116_SLICE_X156Y116_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y116_SLICE_X156Y116_DO5),
.O6(CLBLL_L_X100Y116_SLICE_X156Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff00cc2e2e2e2e)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_CLUT (
.I0(CLBLM_R_X97Y115_SLICE_X153Y115_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y116_SLICE_X160Y116_B5Q),
.I3(CLBLL_L_X100Y116_SLICE_X156Y116_A5Q),
.I4(CLBLL_L_X100Y116_SLICE_X156Y116_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y116_SLICE_X156Y116_CO5),
.O6(CLBLL_L_X100Y116_SLICE_X156Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y116_SLICE_X156Y116_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y116_SLICE_X155Y116_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y116_SLICE_X156Y116_BO5),
.O6(CLBLL_L_X100Y116_SLICE_X156Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X100Y116_SLICE_X156Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y116_SLICE_X156Y116_A5Q),
.I2(CLBLL_L_X100Y117_SLICE_X157Y117_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y116_SLICE_X156Y116_AO5),
.O6(CLBLL_L_X100Y116_SLICE_X156Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X157Y116_AO5),
.Q(CLBLL_L_X100Y116_SLICE_X157Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X157Y116_BO5),
.Q(CLBLL_L_X100Y116_SLICE_X157Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X157Y116_AO6),
.Q(CLBLL_L_X100Y116_SLICE_X157Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y116_SLICE_X157Y116_BO6),
.Q(CLBLL_L_X100Y116_SLICE_X157Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_DLUT (
.I0(CLBLM_L_X98Y115_SLICE_X155Y115_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X100Y116_SLICE_X157Y116_A5Q),
.I4(CLBLL_L_X100Y116_SLICE_X157Y116_AQ),
.I5(CLBLM_R_X97Y115_SLICE_X152Y115_AQ),
.O5(CLBLL_L_X100Y116_SLICE_X157Y116_DO5),
.O6(CLBLL_L_X100Y116_SLICE_X157Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f257f752a207a70)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y117_SLICE_X157Y117_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y118_SLICE_X156Y118_CO6),
.I4(CLBLL_L_X100Y117_SLICE_X157Y117_B5Q),
.I5(CLBLM_L_X92Y116_SLICE_X145Y116_DO6),
.O5(CLBLL_L_X100Y116_SLICE_X157Y116_CO5),
.O6(CLBLL_L_X100Y116_SLICE_X157Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa82828282)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y116_SLICE_X157Y116_A5Q),
.I2(CLBLL_L_X100Y114_SLICE_X156Y114_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X101Y116_SLICE_X158Y116_CO6),
.I5(1'b1),
.O5(CLBLL_L_X100Y116_SLICE_X157Y116_BO5),
.O6(CLBLL_L_X100Y116_SLICE_X157Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLL_L_X100Y116_SLICE_X157Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y116_SLICE_X157Y116_AQ),
.I3(1'b1),
.I4(CLBLM_L_X98Y115_SLICE_X155Y115_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y116_SLICE_X157Y116_AO5),
.O6(CLBLL_L_X100Y116_SLICE_X157Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X156Y117_AO5),
.Q(CLBLL_L_X100Y117_SLICE_X156Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X156Y117_BO5),
.Q(CLBLL_L_X100Y117_SLICE_X156Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X156Y117_AO6),
.Q(CLBLL_L_X100Y117_SLICE_X156Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X156Y117_BO6),
.Q(CLBLL_L_X100Y117_SLICE_X156Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y117_SLICE_X156Y117_AQ),
.I2(CLBLL_L_X100Y117_SLICE_X156Y117_BQ),
.I3(CLBLL_L_X100Y118_SLICE_X156Y118_AQ),
.I4(CLBLL_L_X100Y117_SLICE_X156Y117_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X156Y117_DO5),
.O6(CLBLL_L_X100Y117_SLICE_X156Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f7f43734c7c4070)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_CLUT (
.I0(CLBLL_L_X100Y117_SLICE_X157Y117_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y116_SLICE_X160Y116_C5Q),
.I4(CLBLL_L_X100Y117_SLICE_X156Y117_DO6),
.I5(CLBLM_L_X98Y116_SLICE_X155Y116_DO6),
.O5(CLBLL_L_X100Y117_SLICE_X156Y117_CO5),
.O6(CLBLL_L_X100Y117_SLICE_X156Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y117_SLICE_X156Y117_BQ),
.I2(1'b1),
.I3(CLBLL_L_X100Y118_SLICE_X156Y118_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X156Y117_BO5),
.O6(CLBLL_L_X100Y117_SLICE_X156Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa00aa00aa)
  ) CLBLL_L_X100Y117_SLICE_X156Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X98Y116_SLICE_X155Y116_CO6),
.I4(CLBLL_L_X100Y117_SLICE_X156Y117_CO6),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X156Y117_AO5),
.O6(CLBLL_L_X100Y117_SLICE_X156Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X157Y117_AO5),
.Q(CLBLL_L_X100Y117_SLICE_X157Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X157Y117_BO5),
.Q(CLBLL_L_X100Y117_SLICE_X157Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X157Y117_AO6),
.Q(CLBLL_L_X100Y117_SLICE_X157Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y117_SLICE_X157Y117_BO6),
.Q(CLBLL_L_X100Y117_SLICE_X157Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X157Y117_DO5),
.O6(CLBLL_L_X100Y117_SLICE_X157Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X157Y117_CO5),
.O6(CLBLL_L_X100Y117_SLICE_X157Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y117_SLICE_X158Y117_CO6),
.I2(CLBLM_R_X97Y117_SLICE_X152Y117_BQ),
.I3(CLBLL_L_X100Y118_SLICE_X156Y118_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X157Y117_BO5),
.O6(CLBLL_L_X100Y117_SLICE_X157Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X100Y117_SLICE_X157Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y117_SLICE_X153Y117_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X100Y117_SLICE_X157Y117_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y117_SLICE_X157Y117_AO5),
.O6(CLBLL_L_X100Y117_SLICE_X157Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X156Y118_AO5),
.Q(CLBLL_L_X100Y118_SLICE_X156Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X156Y118_BO5),
.Q(CLBLL_L_X100Y118_SLICE_X156Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X156Y118_AO6),
.Q(CLBLL_L_X100Y118_SLICE_X156Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X156Y118_BO6),
.Q(CLBLL_L_X100Y118_SLICE_X156Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X156Y118_DO5),
.O6(CLBLL_L_X100Y118_SLICE_X156Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_CLUT (
.I0(CLBLL_L_X100Y118_SLICE_X156Y118_BQ),
.I1(CLBLM_L_X92Y116_SLICE_X145Y116_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X100Y118_SLICE_X156Y118_A5Q),
.I4(CLBLL_L_X100Y118_SLICE_X156Y118_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X156Y118_CO5),
.O6(CLBLL_L_X100Y118_SLICE_X156Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y118_SLICE_X156Y118_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y116_SLICE_X145Y116_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X156Y118_BO5),
.O6(CLBLL_L_X100Y118_SLICE_X156Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aa00aa00)
  ) CLBLL_L_X100Y118_SLICE_X156Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X100Y118_SLICE_X156Y118_B5Q),
.I4(CLBLL_L_X100Y117_SLICE_X156Y117_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X156Y118_AO5),
.O6(CLBLL_L_X100Y118_SLICE_X156Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X157Y118_AO5),
.Q(CLBLL_L_X100Y118_SLICE_X157Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X157Y118_BO5),
.Q(CLBLL_L_X100Y118_SLICE_X157Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X157Y118_CO5),
.Q(CLBLL_L_X100Y118_SLICE_X157Y118_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X157Y118_AO6),
.Q(CLBLL_L_X100Y118_SLICE_X157Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X157Y118_BO6),
.Q(CLBLL_L_X100Y118_SLICE_X157Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y118_SLICE_X157Y118_CO6),
.Q(CLBLL_L_X100Y118_SLICE_X157Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X157Y118_DO5),
.O6(CLBLL_L_X100Y118_SLICE_X157Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05050c030c030)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_CLUT (
.I0(CLBLM_R_X103Y117_SLICE_X162Y117_B5Q),
.I1(CLBLL_L_X100Y118_SLICE_X157Y118_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y115_SLICE_X158Y115_A5Q),
.I4(CLBLL_L_X100Y118_SLICE_X157Y118_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X157Y118_CO5),
.O6(CLBLL_L_X100Y118_SLICE_X157Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00aa00a88882222)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y118_SLICE_X157Y118_BQ),
.I2(CLBLM_R_X101Y119_SLICE_X159Y119_B5Q),
.I3(CLBLM_R_X101Y118_SLICE_X158Y118_CQ),
.I4(CLBLL_L_X102Y117_SLICE_X161Y117_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X157Y118_BO5),
.O6(CLBLL_L_X100Y118_SLICE_X157Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLL_L_X100Y118_SLICE_X157Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y119_SLICE_X155Y119_B5Q),
.I2(CLBLL_L_X100Y116_SLICE_X157Y116_B5Q),
.I3(CLBLM_R_X101Y118_SLICE_X159Y118_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y118_SLICE_X157Y118_AO5),
.O6(CLBLL_L_X100Y118_SLICE_X157Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X156Y119_BO5),
.Q(CLBLL_L_X100Y119_SLICE_X156Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X156Y119_AO5),
.Q(CLBLL_L_X100Y119_SLICE_X156Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X156Y119_BO6),
.Q(CLBLL_L_X100Y119_SLICE_X156Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y119_SLICE_X156Y119_DO5),
.O6(CLBLL_L_X100Y119_SLICE_X156Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_CLUT (
.I0(CLBLM_L_X98Y119_SLICE_X155Y119_AQ),
.I1(CLBLL_L_X100Y119_SLICE_X156Y119_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X101Y118_SLICE_X158Y118_CQ),
.I4(CLBLL_L_X100Y119_SLICE_X156Y119_B5Q),
.I5(CLBLM_L_X98Y119_SLICE_X155Y119_BQ),
.O5(CLBLL_L_X100Y119_SLICE_X156Y119_CO5),
.O6(CLBLL_L_X100Y119_SLICE_X156Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y119_SLICE_X155Y119_BQ),
.I2(CLBLL_L_X100Y120_SLICE_X156Y120_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y119_SLICE_X156Y119_BO5),
.O6(CLBLL_L_X100Y119_SLICE_X156Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c88888888)
  ) CLBLL_L_X100Y119_SLICE_X156Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y119_SLICE_X156Y119_B5Q),
.I2(CLBLL_L_X100Y119_SLICE_X156Y119_AQ),
.I3(CLBLM_L_X98Y119_SLICE_X155Y119_BQ),
.I4(CLBLM_L_X98Y119_SLICE_X155Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y119_SLICE_X156Y119_AO5),
.O6(CLBLL_L_X100Y119_SLICE_X156Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X157Y119_BO5),
.Q(CLBLL_L_X100Y119_SLICE_X157Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X157Y119_CO5),
.Q(CLBLL_L_X100Y119_SLICE_X157Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X157Y119_AO6),
.Q(CLBLL_L_X100Y119_SLICE_X157Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y119_SLICE_X157Y119_CO6),
.Q(CLBLL_L_X100Y119_SLICE_X157Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_DLUT (
.I0(CLBLL_L_X100Y119_SLICE_X157Y119_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y120_SLICE_X160Y120_BQ),
.I3(CLBLM_R_X101Y119_SLICE_X158Y119_A5Q),
.I4(CLBLL_L_X100Y119_SLICE_X157Y119_AQ),
.I5(CLBLL_L_X100Y119_SLICE_X157Y119_CQ),
.O5(CLBLL_L_X100Y119_SLICE_X157Y119_DO5),
.O6(CLBLL_L_X100Y119_SLICE_X157Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y119_SLICE_X156Y119_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y119_SLICE_X157Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y119_SLICE_X157Y119_CO5),
.O6(CLBLL_L_X100Y119_SLICE_X157Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c88888888)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y119_SLICE_X158Y119_A5Q),
.I2(CLBLL_L_X100Y119_SLICE_X157Y119_AQ),
.I3(CLBLL_L_X100Y119_SLICE_X157Y119_CQ),
.I4(CLBLL_L_X100Y119_SLICE_X157Y119_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y119_SLICE_X157Y119_BO5),
.O6(CLBLL_L_X100Y119_SLICE_X157Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a8a8202020a820)
  ) CLBLL_L_X100Y119_SLICE_X157Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X92Y120_SLICE_X145Y120_DO6),
.I3(CLBLL_L_X100Y119_SLICE_X157Y119_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y117_SLICE_X155Y117_A5Q),
.O5(CLBLL_L_X100Y119_SLICE_X157Y119_AO5),
.O6(CLBLL_L_X100Y119_SLICE_X157Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y120_SLICE_X156Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y120_SLICE_X156Y120_AO6),
.Q(CLBLL_L_X100Y120_SLICE_X156Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y120_SLICE_X156Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y120_SLICE_X156Y120_DO5),
.O6(CLBLL_L_X100Y120_SLICE_X156Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y120_SLICE_X156Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y120_SLICE_X156Y120_CO5),
.O6(CLBLL_L_X100Y120_SLICE_X156Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y120_SLICE_X156Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y120_SLICE_X156Y120_BO5),
.O6(CLBLL_L_X100Y120_SLICE_X156Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa8a0a8aa0800080)
  ) CLBLL_L_X100Y120_SLICE_X156Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y120_SLICE_X157Y120_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X100Y121_SLICE_X156Y121_AQ),
.I5(CLBLM_L_X92Y119_SLICE_X145Y119_CO6),
.O5(CLBLL_L_X100Y120_SLICE_X156Y120_AO5),
.O6(CLBLL_L_X100Y120_SLICE_X156Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y120_SLICE_X157Y120_AO5),
.Q(CLBLL_L_X100Y120_SLICE_X157Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y120_SLICE_X157Y120_AO6),
.Q(CLBLL_L_X100Y120_SLICE_X157Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y120_SLICE_X157Y120_BO5),
.Q(CLBLL_L_X100Y120_SLICE_X157Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h23202f2ce3e0efec)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_DLUT (
.I0(CLBLM_L_X98Y120_SLICE_X155Y120_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y125_SLICE_X158Y125_CO6),
.I4(CLBLM_R_X97Y120_SLICE_X153Y120_A5Q),
.I5(CLBLL_L_X100Y122_SLICE_X157Y122_BQ),
.O5(CLBLL_L_X100Y120_SLICE_X157Y120_DO5),
.O6(CLBLL_L_X100Y120_SLICE_X157Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_CLUT (
.I0(CLBLL_L_X100Y120_SLICE_X156Y120_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y120_SLICE_X160Y120_B5Q),
.I3(CLBLL_L_X100Y120_SLICE_X157Y120_BQ),
.I4(CLBLL_L_X100Y119_SLICE_X157Y119_C5Q),
.I5(CLBLL_L_X100Y119_SLICE_X156Y119_BQ),
.O5(CLBLL_L_X100Y120_SLICE_X157Y120_CO5),
.O6(CLBLL_L_X100Y120_SLICE_X157Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33ca0a0a0a0)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y120_SLICE_X157Y120_BQ),
.I2(CLBLL_L_X100Y119_SLICE_X157Y119_C5Q),
.I3(CLBLL_L_X100Y119_SLICE_X156Y119_BQ),
.I4(CLBLL_L_X100Y120_SLICE_X156Y120_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y120_SLICE_X157Y120_BO5),
.O6(CLBLL_L_X100Y120_SLICE_X157Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLL_L_X100Y120_SLICE_X157Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y120_SLICE_X157Y120_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y117_SLICE_X155Y117_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y120_SLICE_X157Y120_AO5),
.O6(CLBLL_L_X100Y120_SLICE_X157Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X156Y121_AO5),
.Q(CLBLL_L_X100Y121_SLICE_X156Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X156Y121_CO5),
.Q(CLBLL_L_X100Y121_SLICE_X156Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X156Y121_AO6),
.Q(CLBLL_L_X100Y121_SLICE_X156Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X156Y121_BO6),
.Q(CLBLL_L_X100Y121_SLICE_X156Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X156Y121_CO6),
.Q(CLBLL_L_X100Y121_SLICE_X156Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_DO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_CLUT (
.I0(CLBLM_R_X101Y121_SLICE_X159Y121_C5Q),
.I1(CLBLL_L_X100Y121_SLICE_X156Y121_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y121_SLICE_X159Y121_B5Q),
.I4(CLBLM_R_X97Y121_SLICE_X152Y121_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_CO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa2888022a20080)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLL_L_X100Y121_SLICE_X157Y121_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X93Y121_SLICE_X146Y121_DO6),
.I5(CLBLL_L_X100Y121_SLICE_X156Y121_A5Q),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_BO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y120_SLICE_X157Y120_AQ),
.I3(1'b1),
.I4(CLBLL_L_X100Y121_SLICE_X156Y121_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_AO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X157Y121_CO5),
.Q(CLBLL_L_X100Y121_SLICE_X157Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X157Y121_AO5),
.Q(CLBLL_L_X100Y121_SLICE_X157Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X157Y121_BO6),
.Q(CLBLL_L_X100Y121_SLICE_X157Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y121_SLICE_X157Y121_CO6),
.Q(CLBLL_L_X100Y121_SLICE_X157Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_DLUT (
.I0(CLBLM_L_X98Y121_SLICE_X155Y121_C5Q),
.I1(CLBLL_L_X100Y121_SLICE_X157Y121_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y120_SLICE_X160Y120_DQ),
.I4(CLBLL_L_X100Y121_SLICE_X157Y121_AQ),
.I5(CLBLL_L_X100Y121_SLICE_X156Y121_BQ),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_DO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y120_SLICE_X158Y120_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y121_SLICE_X156Y121_BQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_CO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a82020a820a820)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X93Y121_SLICE_X147Y121_DO6),
.I3(CLBLL_L_X102Y121_SLICE_X160Y121_AO6),
.I4(CLBLL_L_X100Y120_SLICE_X157Y120_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_BO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acccc0000)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_ALUT (
.I0(CLBLL_L_X100Y121_SLICE_X157Y121_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X100Y121_SLICE_X157Y121_AQ),
.I3(CLBLL_L_X100Y121_SLICE_X156Y121_BQ),
.I4(CLBLM_L_X98Y121_SLICE_X155Y121_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_AO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X156Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X156Y122_AO5),
.Q(CLBLL_L_X100Y122_SLICE_X156Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X156Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X156Y122_AO6),
.Q(CLBLL_L_X100Y122_SLICE_X156Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y122_SLICE_X156Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y122_SLICE_X156Y122_DO5),
.O6(CLBLL_L_X100Y122_SLICE_X156Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h73707f7c43404f4c)
  ) CLBLL_L_X100Y122_SLICE_X156Y122_CLUT (
.I0(CLBLM_L_X98Y122_SLICE_X155Y122_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y122_SLICE_X158Y122_DO6),
.I4(CLBLM_R_X97Y121_SLICE_X152Y121_A5Q),
.I5(CLBLM_R_X97Y122_SLICE_X153Y122_DO6),
.O5(CLBLL_L_X100Y122_SLICE_X156Y122_CO5),
.O6(CLBLL_L_X100Y122_SLICE_X156Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111bbbbfa50fa50)
  ) CLBLL_L_X100Y122_SLICE_X156Y122_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y121_SLICE_X156Y121_CQ),
.I2(CLBLM_R_X101Y122_SLICE_X159Y122_DO6),
.I3(CLBLM_R_X101Y121_SLICE_X158Y121_CO6),
.I4(CLBLL_L_X100Y122_SLICE_X156Y122_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X100Y122_SLICE_X156Y122_BO5),
.O6(CLBLL_L_X100Y122_SLICE_X156Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X100Y122_SLICE_X156Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y122_SLICE_X156Y122_A5Q),
.I2(CLBLM_L_X98Y122_SLICE_X155Y122_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y122_SLICE_X156Y122_AO5),
.O6(CLBLL_L_X100Y122_SLICE_X156Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X157Y122_AO5),
.Q(CLBLL_L_X100Y122_SLICE_X157Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X157Y122_BO5),
.Q(CLBLL_L_X100Y122_SLICE_X157Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X157Y122_CO5),
.Q(CLBLL_L_X100Y122_SLICE_X157Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X157Y122_AO6),
.Q(CLBLL_L_X100Y122_SLICE_X157Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X157Y122_BO6),
.Q(CLBLL_L_X100Y122_SLICE_X157Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y122_SLICE_X157Y122_CO6),
.Q(CLBLL_L_X100Y122_SLICE_X157Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y122_SLICE_X157Y122_DO5),
.O6(CLBLL_L_X100Y122_SLICE_X157Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000a0a0a0a0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_CLUT (
.I0(CLBLM_R_X101Y122_SLICE_X158Y122_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y122_SLICE_X157Y122_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y122_SLICE_X157Y122_CO5),
.O6(CLBLL_L_X100Y122_SLICE_X157Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y122_SLICE_X157Y122_CQ),
.I3(CLBLL_L_X100Y122_SLICE_X157Y122_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y122_SLICE_X157Y122_BO5),
.O6(CLBLL_L_X100Y122_SLICE_X157Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030a0a05050)
  ) CLBLL_L_X100Y122_SLICE_X157Y122_ALUT (
.I0(CLBLM_R_X101Y122_SLICE_X159Y122_A5Q),
.I1(CLBLL_L_X100Y122_SLICE_X156Y122_BO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y123_SLICE_X156Y123_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y122_SLICE_X157Y122_AO5),
.O6(CLBLL_L_X100Y122_SLICE_X157Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y123_SLICE_X156Y123_AO5),
.Q(CLBLL_L_X100Y123_SLICE_X156Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y123_SLICE_X156Y123_BO5),
.Q(CLBLL_L_X100Y123_SLICE_X156Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y123_SLICE_X156Y123_AO6),
.Q(CLBLL_L_X100Y123_SLICE_X156Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y123_SLICE_X156Y123_BO6),
.Q(CLBLL_L_X100Y123_SLICE_X156Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_DO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_CO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88228822)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y125_SLICE_X154Y125_A5Q),
.I2(CLBLM_L_X98Y122_SLICE_X155Y122_CO6),
.I3(CLBLM_R_X101Y123_SLICE_X158Y123_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_BO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88228822)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_B5Q),
.I2(CLBLL_L_X100Y122_SLICE_X156Y122_CO6),
.I3(CLBLL_L_X100Y123_SLICE_X156Y123_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_AO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y123_SLICE_X157Y123_AO5),
.Q(CLBLL_L_X100Y123_SLICE_X157Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y123_SLICE_X157Y123_AO6),
.Q(CLBLL_L_X100Y123_SLICE_X157Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_DO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_CO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_BO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y123_SLICE_X157Y123_A5Q),
.I2(CLBLL_L_X100Y122_SLICE_X157Y122_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_AO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X156Y124_BO5),
.Q(CLBLL_L_X100Y124_SLICE_X156Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X156Y124_AO5),
.Q(CLBLL_L_X100Y124_SLICE_X156Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X156Y124_BO6),
.Q(CLBLL_L_X100Y124_SLICE_X156Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y124_SLICE_X156Y124_DO5),
.O6(CLBLL_L_X100Y124_SLICE_X156Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_CLUT (
.I0(CLBLL_L_X100Y124_SLICE_X156Y124_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X98Y125_SLICE_X154Y125_D5Q),
.I3(CLBLL_L_X100Y125_SLICE_X157Y125_DQ),
.I4(CLBLL_L_X100Y124_SLICE_X156Y124_B5Q),
.I5(CLBLL_L_X100Y124_SLICE_X156Y124_AQ),
.O5(CLBLL_L_X100Y124_SLICE_X156Y124_CO5),
.O6(CLBLL_L_X100Y124_SLICE_X156Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaaa0000)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y125_SLICE_X157Y125_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X100Y124_SLICE_X156Y124_BQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y124_SLICE_X156Y124_BO5),
.O6(CLBLL_L_X100Y124_SLICE_X156Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33ca0a0a0a0)
  ) CLBLL_L_X100Y124_SLICE_X156Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y125_SLICE_X157Y125_DQ),
.I2(CLBLL_L_X100Y124_SLICE_X156Y124_B5Q),
.I3(CLBLL_L_X100Y124_SLICE_X156Y124_AQ),
.I4(CLBLL_L_X100Y124_SLICE_X156Y124_BQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y124_SLICE_X156Y124_AO5),
.O6(CLBLL_L_X100Y124_SLICE_X156Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X157Y124_AO5),
.Q(CLBLL_L_X100Y124_SLICE_X157Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X157Y124_BO5),
.Q(CLBLL_L_X100Y124_SLICE_X157Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X157Y124_AO6),
.Q(CLBLL_L_X100Y124_SLICE_X157Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y124_SLICE_X157Y124_BO6),
.Q(CLBLL_L_X100Y124_SLICE_X157Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_DLUT (
.I0(CLBLL_L_X100Y125_SLICE_X157Y125_AQ),
.I1(CLBLL_L_X100Y126_SLICE_X157Y126_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X100Y124_SLICE_X157Y124_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X100Y124_SLICE_X157Y124_AQ),
.O5(CLBLL_L_X100Y124_SLICE_X157Y124_DO5),
.O6(CLBLL_L_X100Y124_SLICE_X157Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22f522a077f577a0)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y123_SLICE_X157Y123_A5Q),
.I2(CLBLM_L_X98Y124_SLICE_X154Y124_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X100Y124_SLICE_X157Y124_DO6),
.I5(CLBLM_R_X97Y121_SLICE_X153Y121_B5Q),
.O5(CLBLL_L_X100Y124_SLICE_X157Y124_CO5),
.O6(CLBLL_L_X100Y124_SLICE_X157Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88882222)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y125_SLICE_X157Y125_C5Q),
.I2(CLBLM_L_X98Y124_SLICE_X154Y124_CO6),
.I3(1'b1),
.I4(CLBLL_L_X100Y124_SLICE_X157Y124_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y124_SLICE_X157Y124_BO5),
.O6(CLBLL_L_X100Y124_SLICE_X157Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLL_L_X100Y124_SLICE_X157Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y124_SLICE_X157Y124_AQ),
.I3(1'b1),
.I4(CLBLL_L_X100Y125_SLICE_X157Y125_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y124_SLICE_X157Y124_AO5),
.O6(CLBLL_L_X100Y124_SLICE_X157Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X156Y125_BO5),
.Q(CLBLL_L_X100Y125_SLICE_X156Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X156Y125_AO6),
.Q(CLBLL_L_X100Y125_SLICE_X156Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X156Y125_BO6),
.Q(CLBLL_L_X100Y125_SLICE_X156Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f1f1f1f0f5f0f5f)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X98Y125_SLICE_X154Y125_C5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X100Y125_SLICE_X156Y125_DO5),
.O6(CLBLL_L_X100Y125_SLICE_X156Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y125_SLICE_X156Y125_AQ),
.I2(CLBLL_L_X100Y125_SLICE_X156Y125_BQ),
.I3(CLBLL_L_X100Y126_SLICE_X156Y126_A5Q),
.I4(CLBLL_L_X100Y125_SLICE_X156Y125_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y125_SLICE_X156Y125_CO5),
.O6(CLBLL_L_X100Y125_SLICE_X156Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y125_SLICE_X156Y125_BQ),
.I2(CLBLL_L_X100Y125_SLICE_X156Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y125_SLICE_X156Y125_BO5),
.O6(CLBLL_L_X100Y125_SLICE_X156Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4055405551555155)
  ) CLBLL_L_X100Y125_SLICE_X156Y125_ALUT (
.I0(CLBLL_L_X100Y125_SLICE_X156Y125_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X100Y126_SLICE_X157Y126_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(1'b1),
.I5(CLBLL_L_X100Y125_SLICE_X156Y125_CO6),
.O5(CLBLL_L_X100Y125_SLICE_X156Y125_AO5),
.O6(CLBLL_L_X100Y125_SLICE_X156Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_AO5),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_BO5),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_CO5),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_AO6),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_BO6),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_CO6),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y125_SLICE_X157Y125_DO6),
.Q(CLBLL_L_X100Y125_SLICE_X157Y125_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa005000d800d800)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y124_SLICE_X156Y124_AO6),
.I2(CLBLL_L_X102Y125_SLICE_X160Y125_DO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X100Y125_SLICE_X157Y125_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X100Y125_SLICE_X157Y125_DO5),
.O6(CLBLL_L_X100Y125_SLICE_X157Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500f0000f00)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_CLUT (
.I0(CLBLL_L_X100Y124_SLICE_X157Y124_CO6),
.I1(1'b1),
.I2(CLBLL_L_X100Y125_SLICE_X157Y125_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X103Y126_SLICE_X163Y126_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y125_SLICE_X157Y125_CO5),
.O6(CLBLL_L_X100Y125_SLICE_X157Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y126_SLICE_X154Y126_AQ),
.I3(CLBLL_L_X100Y125_SLICE_X157Y125_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y125_SLICE_X157Y125_BO5),
.O6(CLBLL_L_X100Y125_SLICE_X157Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X100Y125_SLICE_X157Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y126_SLICE_X157Y126_CQ),
.I2(CLBLM_R_X101Y125_SLICE_X158Y125_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y125_SLICE_X157Y125_AO5),
.O6(CLBLL_L_X100Y125_SLICE_X157Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X156Y126_AO5),
.Q(CLBLL_L_X100Y126_SLICE_X156Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X156Y126_BO5),
.Q(CLBLL_L_X100Y126_SLICE_X156Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X156Y126_AO6),
.Q(CLBLL_L_X100Y126_SLICE_X156Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X156Y126_BO6),
.Q(CLBLL_L_X100Y126_SLICE_X156Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05ff05ff11ff11ff)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLM_L_X98Y126_SLICE_X154Y126_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X100Y126_SLICE_X156Y126_DO5),
.O6(CLBLL_L_X100Y126_SLICE_X156Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y126_SLICE_X156Y126_AQ),
.I2(CLBLL_L_X100Y126_SLICE_X156Y126_BQ),
.I3(1'b1),
.I4(CLBLL_L_X100Y126_SLICE_X156Y126_B5Q),
.I5(CLBLL_L_X100Y126_SLICE_X157Y126_BQ),
.O5(CLBLL_L_X100Y126_SLICE_X156Y126_CO5),
.O6(CLBLL_L_X100Y126_SLICE_X156Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y126_SLICE_X156Y126_BQ),
.I2(CLBLL_L_X100Y126_SLICE_X156Y126_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y126_SLICE_X156Y126_BO5),
.O6(CLBLL_L_X100Y126_SLICE_X156Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000aa00aa00)
  ) CLBLL_L_X100Y126_SLICE_X156Y126_ALUT (
.I0(CLBLL_L_X100Y125_SLICE_X156Y125_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X100Y126_SLICE_X157Y126_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y126_SLICE_X156Y126_AO5),
.O6(CLBLL_L_X100Y126_SLICE_X156Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X157Y126_AO5),
.Q(CLBLL_L_X100Y126_SLICE_X157Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X157Y126_AO6),
.Q(CLBLL_L_X100Y126_SLICE_X157Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X157Y126_BO6),
.Q(CLBLL_L_X100Y126_SLICE_X157Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y126_SLICE_X157Y126_CO6),
.Q(CLBLL_L_X100Y126_SLICE_X157Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055d8d8aaffd8d8)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X98Y127_SLICE_X155Y127_CO6),
.I2(CLBLL_L_X102Y126_SLICE_X160Y126_DO6),
.I3(CLBLM_L_X98Y125_SLICE_X154Y125_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X100Y125_SLICE_X157Y125_BQ),
.O5(CLBLL_L_X100Y126_SLICE_X157Y126_DO5),
.O6(CLBLL_L_X100Y126_SLICE_X157Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3131333311111313)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y126_SLICE_X158Y126_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y124_SLICE_X157Y124_DO6),
.I5(CLBLM_R_X101Y126_SLICE_X158Y126_AQ),
.O5(CLBLL_L_X100Y126_SLICE_X157Y126_CO5),
.O6(CLBLL_L_X100Y126_SLICE_X157Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h008b00ff008b00ff)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_BLUT (
.I0(CLBLL_L_X100Y126_SLICE_X157Y126_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X100Y126_SLICE_X156Y126_CO6),
.I3(CLBLL_L_X100Y126_SLICE_X156Y126_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLL_L_X100Y126_SLICE_X157Y126_BO5),
.O6(CLBLL_L_X100Y126_SLICE_X157Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLL_L_X100Y126_SLICE_X157Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y126_SLICE_X157Y126_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X101Y126_SLICE_X158Y126_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y126_SLICE_X157Y126_AO5),
.O6(CLBLL_L_X100Y126_SLICE_X157Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X156Y127_AO5),
.Q(CLBLL_L_X100Y127_SLICE_X156Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X156Y127_BO5),
.Q(CLBLL_L_X100Y127_SLICE_X156Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X156Y127_AO6),
.Q(CLBLL_L_X100Y127_SLICE_X156Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X156Y127_BO6),
.Q(CLBLL_L_X100Y127_SLICE_X156Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y127_SLICE_X156Y127_DO5),
.O6(CLBLL_L_X100Y127_SLICE_X156Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y127_SLICE_X156Y127_BQ),
.I3(CLBLL_L_X100Y127_SLICE_X156Y127_A5Q),
.I4(CLBLL_L_X100Y127_SLICE_X156Y127_B5Q),
.I5(CLBLL_L_X100Y128_SLICE_X156Y128_BQ),
.O5(CLBLL_L_X100Y127_SLICE_X156Y127_CO5),
.O6(CLBLL_L_X100Y127_SLICE_X156Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X100Y128_SLICE_X156Y128_BQ),
.I4(CLBLL_L_X100Y127_SLICE_X156Y127_BQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y127_SLICE_X156Y127_BO5),
.O6(CLBLL_L_X100Y127_SLICE_X156Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLL_L_X100Y127_SLICE_X156Y127_ALUT (
.I0(CLBLL_L_X100Y127_SLICE_X156Y127_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X100Y127_SLICE_X157Y127_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y127_SLICE_X156Y127_AO5),
.O6(CLBLL_L_X100Y127_SLICE_X156Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X157Y127_BO5),
.Q(CLBLL_L_X100Y127_SLICE_X157Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X157Y127_AO6),
.Q(CLBLL_L_X100Y127_SLICE_X157Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y127_SLICE_X157Y127_BO6),
.Q(CLBLL_L_X100Y127_SLICE_X157Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y127_SLICE_X157Y127_DO5),
.O6(CLBLL_L_X100Y127_SLICE_X157Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_CLUT (
.I0(CLBLL_L_X100Y127_SLICE_X156Y127_AQ),
.I1(1'b1),
.I2(CLBLL_L_X100Y127_SLICE_X157Y127_BQ),
.I3(CLBLL_L_X100Y127_SLICE_X157Y127_AQ),
.I4(CLBLL_L_X100Y127_SLICE_X157Y127_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X100Y127_SLICE_X157Y127_CO5),
.O6(CLBLL_L_X100Y127_SLICE_X157Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y127_SLICE_X157Y127_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X100Y127_SLICE_X156Y127_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y127_SLICE_X157Y127_BO5),
.O6(CLBLL_L_X100Y127_SLICE_X157Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2323030333331313)
  ) CLBLL_L_X100Y127_SLICE_X157Y127_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X100Y129_SLICE_X157Y129_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y128_SLICE_X156Y128_AQ),
.I5(CLBLL_L_X100Y127_SLICE_X157Y127_CO6),
.O5(CLBLL_L_X100Y127_SLICE_X157Y127_AO5),
.O6(CLBLL_L_X100Y127_SLICE_X157Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y128_SLICE_X156Y128_AO5),
.Q(CLBLL_L_X100Y128_SLICE_X156Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y128_SLICE_X156Y128_AO6),
.Q(CLBLL_L_X100Y128_SLICE_X156Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y128_SLICE_X156Y128_BO6),
.Q(CLBLL_L_X100Y128_SLICE_X156Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y128_SLICE_X156Y128_DO5),
.O6(CLBLL_L_X100Y128_SLICE_X156Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555557777557777)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_L_X98Y127_SLICE_X154Y127_B5Q),
.O5(CLBLL_L_X100Y128_SLICE_X156Y128_CO5),
.O6(CLBLL_L_X100Y128_SLICE_X156Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff3f0f3f)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y127_SLICE_X156Y127_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X100Y128_SLICE_X156Y128_A5Q),
.I5(CLBLL_L_X100Y128_SLICE_X156Y128_CO6),
.O5(CLBLL_L_X100Y128_SLICE_X156Y128_BO5),
.O6(CLBLL_L_X100Y128_SLICE_X156Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLL_L_X100Y128_SLICE_X156Y128_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y128_SLICE_X156Y128_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y126_SLICE_X157Y126_AQ),
.I5(1'b1),
.O5(CLBLL_L_X100Y128_SLICE_X156Y128_AO5),
.O6(CLBLL_L_X100Y128_SLICE_X156Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y128_SLICE_X157Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y128_SLICE_X157Y128_DO5),
.O6(CLBLL_L_X100Y128_SLICE_X157Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y128_SLICE_X157Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y128_SLICE_X157Y128_CO5),
.O6(CLBLL_L_X100Y128_SLICE_X157Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y128_SLICE_X157Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y128_SLICE_X157Y128_BO5),
.O6(CLBLL_L_X100Y128_SLICE_X157Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y128_SLICE_X157Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y128_SLICE_X157Y128_AO5),
.O6(CLBLL_L_X100Y128_SLICE_X157Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y129_SLICE_X156Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y129_SLICE_X156Y129_AO6),
.Q(CLBLL_L_X100Y129_SLICE_X156Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y129_SLICE_X156Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y129_SLICE_X156Y129_DO5),
.O6(CLBLL_L_X100Y129_SLICE_X156Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y129_SLICE_X156Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y129_SLICE_X156Y129_CO5),
.O6(CLBLL_L_X100Y129_SLICE_X156Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5752f7f20702a7a2)
  ) CLBLL_L_X100Y129_SLICE_X156Y129_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X98Y128_SLICE_X154Y128_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y129_SLICE_X158Y129_CO6),
.I4(CLBLM_L_X98Y129_SLICE_X155Y129_AQ),
.I5(CLBLM_L_X98Y128_SLICE_X154Y128_DO6),
.O5(CLBLL_L_X100Y129_SLICE_X156Y129_BO5),
.O6(CLBLL_L_X100Y129_SLICE_X156Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cc00cc0c00cc00c)
  ) CLBLL_L_X100Y129_SLICE_X156Y129_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X100Y130_SLICE_X156Y130_AQ),
.I3(CLBLM_L_X98Y128_SLICE_X154Y128_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X97Y128_SLICE_X153Y128_A5Q),
.O5(CLBLL_L_X100Y129_SLICE_X156Y129_AO5),
.O6(CLBLL_L_X100Y129_SLICE_X156Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y129_SLICE_X157Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y129_SLICE_X157Y129_AO5),
.Q(CLBLL_L_X100Y129_SLICE_X157Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y129_SLICE_X157Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y129_SLICE_X157Y129_AO6),
.Q(CLBLL_L_X100Y129_SLICE_X157Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y129_SLICE_X157Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y129_SLICE_X157Y129_DO5),
.O6(CLBLL_L_X100Y129_SLICE_X157Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y129_SLICE_X157Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y129_SLICE_X157Y129_CO5),
.O6(CLBLL_L_X100Y129_SLICE_X157Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0505ffffffff)
  ) CLBLL_L_X100Y129_SLICE_X157Y129_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y127_SLICE_X155Y127_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLL_L_X100Y129_SLICE_X157Y129_BO5),
.O6(CLBLL_L_X100Y129_SLICE_X157Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLL_L_X100Y129_SLICE_X157Y129_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y129_SLICE_X156Y129_BO6),
.I2(CLBLM_L_X98Y127_SLICE_X155Y127_A5Q),
.I3(CLBLM_R_X101Y130_SLICE_X158Y130_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y129_SLICE_X157Y129_AO5),
.O6(CLBLL_L_X100Y129_SLICE_X157Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y130_SLICE_X156Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y130_SLICE_X156Y130_AO6),
.Q(CLBLL_L_X100Y130_SLICE_X156Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X156Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X156Y130_DO5),
.O6(CLBLL_L_X100Y130_SLICE_X156Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X156Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X156Y130_CO5),
.O6(CLBLL_L_X100Y130_SLICE_X156Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X156Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X156Y130_BO5),
.O6(CLBLL_L_X100Y130_SLICE_X156Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0055005500)
  ) CLBLL_L_X100Y130_SLICE_X156Y130_ALUT (
.I0(CLBLL_L_X100Y133_SLICE_X156Y133_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(CLBLM_L_X98Y130_SLICE_X154Y130_A5Q),
.O5(CLBLL_L_X100Y130_SLICE_X156Y130_AO5),
.O6(CLBLL_L_X100Y130_SLICE_X156Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X157Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X157Y130_DO5),
.O6(CLBLL_L_X100Y130_SLICE_X157Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X157Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X157Y130_CO5),
.O6(CLBLL_L_X100Y130_SLICE_X157Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X157Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X157Y130_BO5),
.O6(CLBLL_L_X100Y130_SLICE_X157Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y130_SLICE_X157Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y130_SLICE_X157Y130_AO5),
.O6(CLBLL_L_X100Y130_SLICE_X157Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y133_SLICE_X156Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y133_SLICE_X156Y133_AO5),
.Q(CLBLL_L_X100Y133_SLICE_X156Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y133_SLICE_X156Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y133_SLICE_X156Y133_AO6),
.Q(CLBLL_L_X100Y133_SLICE_X156Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X156Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X156Y133_DO5),
.O6(CLBLL_L_X100Y133_SLICE_X156Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X156Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X156Y133_CO5),
.O6(CLBLL_L_X100Y133_SLICE_X156Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X156Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X156Y133_BO5),
.O6(CLBLL_L_X100Y133_SLICE_X156Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0000aa82828282)
  ) CLBLL_L_X100Y133_SLICE_X156Y133_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y133_SLICE_X152Y133_A5Q),
.I2(CLBLL_L_X100Y133_SLICE_X156Y133_AQ),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_A5Q),
.I4(CLBLL_L_X100Y134_SLICE_X156Y134_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X156Y133_AO5),
.O6(CLBLL_L_X100Y133_SLICE_X156Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X157Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X157Y133_DO5),
.O6(CLBLL_L_X100Y133_SLICE_X157Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X157Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X157Y133_CO5),
.O6(CLBLL_L_X100Y133_SLICE_X157Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X157Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X157Y133_BO5),
.O6(CLBLL_L_X100Y133_SLICE_X157Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y133_SLICE_X157Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y133_SLICE_X157Y133_AO5),
.O6(CLBLL_L_X100Y133_SLICE_X157Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y134_SLICE_X156Y134_AO5),
.Q(CLBLL_L_X100Y134_SLICE_X156Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y134_SLICE_X156Y134_BO5),
.Q(CLBLL_L_X100Y134_SLICE_X156Y134_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y134_SLICE_X156Y134_AO6),
.Q(CLBLL_L_X100Y134_SLICE_X156Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X100Y134_SLICE_X156Y134_BO6),
.Q(CLBLL_L_X100Y134_SLICE_X156Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X156Y134_DO5),
.O6(CLBLL_L_X100Y134_SLICE_X156Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3cc3aaaac33c)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_CLUT (
.I0(CLBLM_L_X98Y132_SLICE_X155Y132_C5Q),
.I1(CLBLM_R_X101Y134_SLICE_X158Y134_AQ),
.I2(CLBLL_L_X100Y134_SLICE_X156Y134_AQ),
.I3(CLBLL_L_X100Y134_SLICE_X156Y134_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X101Y134_SLICE_X159Y134_BQ),
.O5(CLBLL_L_X100Y134_SLICE_X156Y134_CO5),
.O6(CLBLL_L_X100Y134_SLICE_X156Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa005500c300c300)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_BLUT (
.I0(CLBLM_R_X97Y133_SLICE_X153Y133_A5Q),
.I1(CLBLL_L_X100Y134_SLICE_X156Y134_BQ),
.I2(CLBLM_L_X98Y134_SLICE_X154Y134_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y132_SLICE_X155Y132_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X156Y134_BO5),
.O6(CLBLL_L_X100Y134_SLICE_X156Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLL_L_X100Y134_SLICE_X156Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y134_SLICE_X158Y134_AQ),
.I2(CLBLL_L_X100Y134_SLICE_X156Y134_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X156Y134_AO5),
.O6(CLBLL_L_X100Y134_SLICE_X156Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y134_SLICE_X157Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X157Y134_DO5),
.O6(CLBLL_L_X100Y134_SLICE_X157Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y134_SLICE_X157Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X157Y134_CO5),
.O6(CLBLL_L_X100Y134_SLICE_X157Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y134_SLICE_X157Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X157Y134_BO5),
.O6(CLBLL_L_X100Y134_SLICE_X157Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y134_SLICE_X157Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y134_SLICE_X157Y134_AO5),
.O6(CLBLL_L_X100Y134_SLICE_X157Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_BO5),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_BO6),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y112_SLICE_X159Y112_C5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y111_SLICE_X160Y111_BQ),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q),
.I5(CLBLM_R_X101Y112_SLICE_X158Y112_BQ),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_DO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h47474747ffcc3300)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_CLUT (
.I0(CLBLL_L_X102Y111_SLICE_X161Y111_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLL_L_X102Y111_SLICE_X161Y111_B5Q),
.I3(CLBLM_R_X101Y112_SLICE_X158Y112_CO6),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_CO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y111_SLICE_X160Y111_BQ),
.I2(1'b1),
.I3(CLBLM_R_X101Y112_SLICE_X158Y112_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_BO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f00ffaaaa0000)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y111_SLICE_X160Y111_DO6),
.I4(CLBLL_L_X102Y111_SLICE_X161Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_AO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y111_SLICE_X161Y111_BO5),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y111_SLICE_X161Y111_AO5),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y111_SLICE_X161Y111_BO6),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_AO5),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff0fcc55000fcc)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_DLUT (
.I0(CLBLM_R_X103Y111_SLICE_X162Y111_AQ),
.I1(CLBLM_R_X101Y111_SLICE_X158Y111_DO6),
.I2(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X103Y111_SLICE_X162Y111_CO6),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_DO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30773044fc77fc44)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_CLUT (
.I0(CLBLL_L_X102Y111_SLICE_X161Y111_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y112_SLICE_X162Y112_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLL_L_X100Y111_SLICE_X156Y111_DO6),
.I5(CLBLL_L_X102Y111_SLICE_X161Y111_CQ),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_CO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00a0a88228822)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y111_SLICE_X161Y111_BQ),
.I2(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q),
.I3(CLBLM_R_X101Y112_SLICE_X159Y112_C5Q),
.I4(CLBLM_R_X103Y112_SLICE_X162Y112_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_BO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc03fc03fa0a0a0a0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y111_SLICE_X161Y111_CQ),
.I3(CLBLM_R_X103Y112_SLICE_X162Y112_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_AO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_BO5),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_AO5),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_BO6),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_AO5),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_DLUT (
.I0(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I1(1'b1),
.I2(CLBLL_L_X100Y112_SLICE_X157Y112_AQ),
.I3(CLBLM_R_X101Y112_SLICE_X159Y112_CQ),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_DO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f5f5030305f50)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_CLUT (
.I0(CLBLL_L_X102Y113_SLICE_X160Y113_AQ),
.I1(CLBLL_L_X102Y112_SLICE_X160Y112_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y112_SLICE_X156Y112_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y112_SLICE_X160Y112_DO6),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_CO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaaa0000)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y112_SLICE_X159Y112_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_BO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc03fc03fa0a0a0a0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_CQ),
.I3(CLBLL_L_X102Y112_SLICE_X160Y112_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_AO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_AO5),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_BO5),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_AO6),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_BO6),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_DO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505fcfcf505fc0c0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_CLUT (
.I0(CLBLM_R_X103Y112_SLICE_X163Y112_BQ),
.I1(CLBLM_R_X103Y112_SLICE_X163Y112_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X101Y110_SLICE_X158Y110_CO6),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_CO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00aa00a88882222)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I2(CLBLL_L_X102Y113_SLICE_X161Y113_B5Q),
.I3(CLBLM_R_X103Y112_SLICE_X163Y112_A5Q),
.I4(CLBLM_R_X103Y112_SLICE_X162Y112_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_BO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y113_SLICE_X161Y113_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X101Y110_SLICE_X158Y110_A5Q),
.I4(CLBLL_L_X102Y112_SLICE_X161Y112_CO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_AO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y113_SLICE_X160Y113_AO5),
.Q(CLBLL_L_X102Y113_SLICE_X160Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y113_SLICE_X160Y113_AO6),
.Q(CLBLL_L_X102Y113_SLICE_X160Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_DO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_CO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_BO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa550000c3c30000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_ALUT (
.I0(CLBLL_L_X102Y111_SLICE_X161Y111_B5Q),
.I1(CLBLM_R_X101Y113_SLICE_X158Y113_A5Q),
.I2(CLBLL_L_X102Y113_SLICE_X160Y113_AQ),
.I3(CLBLL_L_X102Y112_SLICE_X160Y112_B5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_AO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y113_SLICE_X161Y113_AO5),
.Q(CLBLL_L_X102Y113_SLICE_X161Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y113_SLICE_X161Y113_BO5),
.Q(CLBLL_L_X102Y113_SLICE_X161Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y113_SLICE_X161Y113_AO6),
.Q(CLBLL_L_X102Y113_SLICE_X161Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y113_SLICE_X161Y113_BO6),
.Q(CLBLL_L_X102Y113_SLICE_X161Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h505ffcfc505f0c0c)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_DLUT (
.I0(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I1(CLBLM_R_X101Y113_SLICE_X159Y113_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X102Y113_SLICE_X161Y113_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X102Y114_SLICE_X161Y114_BO6),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_DO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ca0fcaf0caffca)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_CLUT (
.I0(CLBLM_R_X101Y112_SLICE_X159Y112_DO6),
.I1(CLBLM_R_X103Y113_SLICE_X162Y113_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y113_SLICE_X161Y113_B5Q),
.I5(CLBLM_R_X103Y113_SLICE_X163Y113_AQ),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_CO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00a0a88228822)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y113_SLICE_X161Y113_BQ),
.I2(CLBLL_L_X102Y114_SLICE_X161Y114_A5Q),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q),
.I4(CLBLL_L_X102Y115_SLICE_X161Y115_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_BO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa82828282)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y112_SLICE_X159Y112_B5Q),
.I2(CLBLL_L_X102Y114_SLICE_X160Y114_B5Q),
.I3(1'b1),
.I4(CLBLL_L_X102Y113_SLICE_X161Y113_CO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_AO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X160Y114_BO5),
.Q(CLBLL_L_X102Y114_SLICE_X160Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X160Y114_CO5),
.Q(CLBLL_L_X102Y114_SLICE_X160Y114_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X160Y114_BO6),
.Q(CLBLL_L_X102Y114_SLICE_X160Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X160Y114_CO6),
.Q(CLBLL_L_X102Y114_SLICE_X160Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_DO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cc00cc00)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X102Y114_SLICE_X160Y114_BQ),
.I3(CLBLL_L_X102Y115_SLICE_X160Y115_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_CO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc84848484)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_BLUT (
.I0(CLBLL_L_X102Y115_SLICE_X160Y115_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y112_SLICE_X159Y112_A5Q),
.I3(CLBLL_L_X102Y113_SLICE_X161Y113_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_BO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0055ffcc00cc00)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X102Y115_SLICE_X160Y115_CQ),
.I4(CLBLL_L_X102Y115_SLICE_X160Y115_DO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_AO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X161Y114_AO5),
.Q(CLBLL_L_X102Y114_SLICE_X161Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X161Y114_AO6),
.Q(CLBLL_L_X102Y114_SLICE_X161Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_DO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_CO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y114_SLICE_X160Y114_CQ),
.I2(CLBLL_L_X102Y114_SLICE_X161Y114_AQ),
.I3(CLBLL_L_X102Y114_SLICE_X160Y114_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y114_SLICE_X161Y114_A5Q),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_BO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y114_SLICE_X160Y114_CQ),
.I2(CLBLL_L_X102Y114_SLICE_X161Y114_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_AO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X160Y115_AO5),
.Q(CLBLL_L_X102Y115_SLICE_X160Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X160Y115_BO5),
.Q(CLBLL_L_X102Y115_SLICE_X160Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X160Y115_AO6),
.Q(CLBLL_L_X102Y115_SLICE_X160Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X160Y115_BO6),
.Q(CLBLL_L_X102Y115_SLICE_X160Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_AO5),
.Q(CLBLL_L_X102Y115_SLICE_X160Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_DLUT (
.I0(CLBLL_L_X102Y114_SLICE_X160Y114_C5Q),
.I1(CLBLL_L_X102Y115_SLICE_X160Y115_AQ),
.I2(CLBLL_L_X102Y115_SLICE_X160Y115_BQ),
.I3(1'b1),
.I4(CLBLL_L_X102Y115_SLICE_X160Y115_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_DO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22fa225077fa7750)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y115_SLICE_X160Y115_CQ),
.I2(CLBLM_R_X101Y116_SLICE_X158Y116_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y115_SLICE_X160Y115_DO6),
.I5(CLBLL_L_X102Y115_SLICE_X161Y115_C5Q),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_CO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X102Y115_SLICE_X160Y115_AQ),
.I3(1'b1),
.I4(CLBLL_L_X102Y115_SLICE_X160Y115_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_BO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00a500a500)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_ALUT (
.I0(CLBLM_R_X101Y116_SLICE_X158Y116_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X102Y116_SLICE_X160Y116_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y115_SLICE_X160Y115_CO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_AO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_BO5),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_CO5),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_BO6),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_CO6),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y116_SLICE_X160Y116_CQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_BQ),
.I4(CLBLL_L_X102Y115_SLICE_X161Y115_B5Q),
.I5(CLBLL_L_X102Y116_SLICE_X161Y116_A5Q),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_DO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_CLUT (
.I0(CLBLL_L_X102Y114_SLICE_X160Y114_C5Q),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y117_SLICE_X158Y117_B5Q),
.I4(CLBLL_L_X102Y116_SLICE_X161Y116_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_CO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_BLUT (
.I0(CLBLL_L_X102Y116_SLICE_X160Y116_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y115_SLICE_X161Y115_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_BO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5500ffcccc0000)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X102Y116_SLICE_X161Y116_DO6),
.I4(CLBLL_L_X102Y116_SLICE_X161Y116_CQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_AO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X160Y116_BO5),
.Q(CLBLL_L_X102Y116_SLICE_X160Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X160Y116_CO5),
.Q(CLBLL_L_X102Y116_SLICE_X160Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X159Y116_AO5),
.Q(CLBLL_L_X102Y116_SLICE_X160Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X160Y116_BO6),
.Q(CLBLL_L_X102Y116_SLICE_X160Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X160Y116_CO6),
.Q(CLBLL_L_X102Y116_SLICE_X160Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2727ff552727aa00)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y116_SLICE_X160Y116_AQ),
.I2(CLBLM_R_X101Y117_SLICE_X158Y117_B5Q),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X100Y117_SLICE_X156Y117_DO6),
.O5(CLBLL_L_X102Y116_SLICE_X160Y116_DO5),
.O6(CLBLL_L_X102Y116_SLICE_X160Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00c300c300)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y117_SLICE_X156Y117_B5Q),
.I2(CLBLL_L_X100Y117_SLICE_X157Y117_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y116_SLICE_X160Y116_DO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y116_SLICE_X160Y116_CO5),
.O6(CLBLL_L_X102Y116_SLICE_X160Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00aa005500)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_BLUT (
.I0(CLBLM_R_X101Y116_SLICE_X158Y116_A5Q),
.I1(1'b1),
.I2(CLBLL_L_X102Y116_SLICE_X161Y116_CO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y116_SLICE_X160Y116_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y116_SLICE_X160Y116_BO5),
.O6(CLBLL_L_X102Y116_SLICE_X160Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05fc0c0c0c0)
  ) CLBLL_L_X102Y116_SLICE_X160Y116_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X102Y116_SLICE_X160Y116_AQ),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y116_SLICE_X160Y116_AO5),
.O6(CLBLL_L_X102Y116_SLICE_X160Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X161Y116_AO5),
.Q(CLBLL_L_X102Y116_SLICE_X161Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X161Y116_BO5),
.Q(CLBLL_L_X102Y116_SLICE_X161Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X161Y116_AO6),
.Q(CLBLL_L_X102Y116_SLICE_X161Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X161Y116_BO6),
.Q(CLBLL_L_X102Y116_SLICE_X161Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y116_SLICE_X160Y116_AO5),
.Q(CLBLL_L_X102Y116_SLICE_X161Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y116_SLICE_X161Y116_AQ),
.I2(CLBLL_L_X102Y116_SLICE_X161Y116_BQ),
.I3(1'b1),
.I4(CLBLL_L_X102Y116_SLICE_X161Y116_B5Q),
.I5(CLBLL_L_X102Y116_SLICE_X160Y116_BQ),
.O5(CLBLL_L_X102Y116_SLICE_X161Y116_DO5),
.O6(CLBLL_L_X102Y116_SLICE_X161Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22772277fafa5050)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y116_SLICE_X161Y116_CQ),
.I2(CLBLL_L_X100Y116_SLICE_X156Y116_DO6),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_CQ),
.I4(CLBLL_L_X102Y116_SLICE_X161Y116_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y116_SLICE_X161Y116_CO5),
.O6(CLBLL_L_X102Y116_SLICE_X161Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y116_SLICE_X161Y116_BQ),
.I2(CLBLL_L_X102Y116_SLICE_X161Y116_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y116_SLICE_X161Y116_BO5),
.O6(CLBLL_L_X102Y116_SLICE_X161Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLL_L_X102Y116_SLICE_X161Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_B5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y116_SLICE_X160Y116_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y116_SLICE_X161Y116_AO5),
.O6(CLBLL_L_X102Y116_SLICE_X161Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X160Y117_BO5),
.Q(CLBLL_L_X102Y117_SLICE_X160Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X160Y117_AO6),
.Q(CLBLL_L_X102Y117_SLICE_X160Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X160Y117_BO6),
.Q(CLBLL_L_X102Y117_SLICE_X160Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699696696996)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_DLUT (
.I0(CLBLM_R_X101Y117_SLICE_X159Y117_BQ),
.I1(CLBLL_L_X102Y117_SLICE_X160Y117_AQ),
.I2(CLBLL_L_X102Y117_SLICE_X160Y117_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y117_SLICE_X160Y117_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y117_SLICE_X160Y117_DO5),
.O6(CLBLL_L_X102Y117_SLICE_X160Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996696696996)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_CLUT (
.I0(CLBLM_R_X101Y117_SLICE_X159Y117_BQ),
.I1(CLBLL_L_X102Y117_SLICE_X160Y117_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y117_SLICE_X160Y117_BQ),
.I4(CLBLL_L_X102Y117_SLICE_X160Y117_B5Q),
.I5(CLBLL_L_X102Y117_SLICE_X161Y117_C5Q),
.O5(CLBLL_L_X102Y117_SLICE_X160Y117_CO5),
.O6(CLBLL_L_X102Y117_SLICE_X160Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_BLUT (
.I0(CLBLL_L_X102Y117_SLICE_X160Y117_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y117_SLICE_X159Y117_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y117_SLICE_X160Y117_BO5),
.O6(CLBLL_L_X102Y117_SLICE_X160Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he200ff00e2000000)
  ) CLBLL_L_X102Y117_SLICE_X160Y117_ALUT (
.I0(CLBLL_L_X102Y117_SLICE_X160Y117_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y117_SLICE_X161Y117_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X100Y119_SLICE_X156Y119_CO6),
.O5(CLBLL_L_X102Y117_SLICE_X160Y117_AO5),
.O6(CLBLL_L_X102Y117_SLICE_X160Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_AO5),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_BO5),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_CO5),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_DO5),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_AO6),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_BO6),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_CO6),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y117_SLICE_X161Y117_DO6),
.Q(CLBLL_L_X102Y117_SLICE_X161Y117_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y117_SLICE_X162Y117_AQ),
.I3(CLBLM_R_X103Y116_SLICE_X162Y116_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y117_SLICE_X161Y117_DO5),
.O6(CLBLL_L_X102Y117_SLICE_X161Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y122_SLICE_X160Y122_BQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y117_SLICE_X161Y117_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y117_SLICE_X161Y117_CO5),
.O6(CLBLL_L_X102Y117_SLICE_X161Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888c0c0c0c0)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_BLUT (
.I0(CLBLL_L_X102Y117_SLICE_X161Y117_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X102Y117_SLICE_X161Y117_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y117_SLICE_X161Y117_BO5),
.O6(CLBLL_L_X102Y117_SLICE_X161Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLL_L_X102Y117_SLICE_X161Y117_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y117_SLICE_X161Y117_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y117_SLICE_X161Y117_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y117_SLICE_X161Y117_AO5),
.O6(CLBLL_L_X102Y117_SLICE_X161Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X160Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X160Y118_DO5),
.O6(CLBLL_L_X102Y118_SLICE_X160Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X160Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X160Y118_CO5),
.O6(CLBLL_L_X102Y118_SLICE_X160Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X160Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X160Y118_BO5),
.O6(CLBLL_L_X102Y118_SLICE_X160Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c03f3f22222222)
  ) CLBLL_L_X102Y118_SLICE_X160Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y118_SLICE_X159Y118_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(1'b1),
.I4(CLBLM_R_X101Y118_SLICE_X159Y118_DO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X160Y118_AO5),
.O6(CLBLL_L_X102Y118_SLICE_X160Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X161Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X161Y118_DO5),
.O6(CLBLL_L_X102Y118_SLICE_X161Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X161Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X161Y118_CO5),
.O6(CLBLL_L_X102Y118_SLICE_X161Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X161Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X161Y118_BO5),
.O6(CLBLL_L_X102Y118_SLICE_X161Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y118_SLICE_X161Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y118_SLICE_X161Y118_AO5),
.O6(CLBLL_L_X102Y118_SLICE_X161Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X160Y119_AO5),
.Q(CLBLL_L_X102Y119_SLICE_X160Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X160Y119_BO5),
.Q(CLBLL_L_X102Y119_SLICE_X160Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X160Y119_AO6),
.Q(CLBLL_L_X102Y119_SLICE_X160Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X160Y119_BO6),
.Q(CLBLL_L_X102Y119_SLICE_X160Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696696969699696)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_DLUT (
.I0(CLBLL_L_X102Y120_SLICE_X160Y120_AQ),
.I1(CLBLL_L_X102Y119_SLICE_X160Y119_AQ),
.I2(CLBLL_L_X102Y119_SLICE_X160Y119_BQ),
.I3(1'b1),
.I4(CLBLL_L_X102Y119_SLICE_X160Y119_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y119_SLICE_X160Y119_DO5),
.O6(CLBLL_L_X102Y119_SLICE_X160Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h699696695aa5a55a)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_CLUT (
.I0(CLBLL_L_X102Y120_SLICE_X160Y120_AQ),
.I1(CLBLM_R_X103Y120_SLICE_X162Y120_CQ),
.I2(CLBLL_L_X102Y119_SLICE_X160Y119_AQ),
.I3(CLBLL_L_X102Y119_SLICE_X160Y119_BQ),
.I4(CLBLL_L_X102Y119_SLICE_X160Y119_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y119_SLICE_X160Y119_CO5),
.O6(CLBLL_L_X102Y119_SLICE_X160Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y119_SLICE_X160Y119_BQ),
.I2(CLBLL_L_X102Y119_SLICE_X160Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y119_SLICE_X160Y119_BO5),
.O6(CLBLL_L_X102Y119_SLICE_X160Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X102Y119_SLICE_X160Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y119_SLICE_X161Y119_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y120_SLICE_X160Y120_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y119_SLICE_X160Y119_AO5),
.O6(CLBLL_L_X102Y119_SLICE_X160Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X161Y119_BO5),
.Q(CLBLL_L_X102Y119_SLICE_X161Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X161Y119_AO6),
.Q(CLBLL_L_X102Y119_SLICE_X161Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y119_SLICE_X161Y119_BO6),
.Q(CLBLL_L_X102Y119_SLICE_X161Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966669966999966)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_DLUT (
.I0(CLBLL_L_X102Y119_SLICE_X161Y119_BQ),
.I1(CLBLL_L_X102Y119_SLICE_X160Y119_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y119_SLICE_X161Y119_B5Q),
.I5(CLBLL_L_X102Y119_SLICE_X161Y119_AQ),
.O5(CLBLL_L_X102Y119_SLICE_X161Y119_DO5),
.O6(CLBLL_L_X102Y119_SLICE_X161Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966969996996966)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_CLUT (
.I0(CLBLL_L_X102Y119_SLICE_X161Y119_BQ),
.I1(CLBLL_L_X102Y119_SLICE_X160Y119_A5Q),
.I2(CLBLM_R_X103Y120_SLICE_X162Y120_C5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y119_SLICE_X161Y119_B5Q),
.I5(CLBLL_L_X102Y119_SLICE_X161Y119_AQ),
.O5(CLBLL_L_X102Y119_SLICE_X161Y119_CO5),
.O6(CLBLL_L_X102Y119_SLICE_X161Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y119_SLICE_X161Y119_BQ),
.I2(CLBLL_L_X102Y119_SLICE_X161Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y119_SLICE_X161Y119_BO5),
.O6(CLBLL_L_X102Y119_SLICE_X161Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa00a0088888888)
  ) CLBLL_L_X102Y119_SLICE_X161Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y120_SLICE_X158Y120_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y119_SLICE_X161Y119_DO6),
.I4(CLBLM_R_X103Y120_SLICE_X162Y120_C5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLL_L_X102Y119_SLICE_X161Y119_AO5),
.O6(CLBLL_L_X102Y119_SLICE_X161Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_BO5),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_CO5),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_DO5),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_AO6),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_BO6),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_CO6),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X160Y120_DO6),
.Q(CLBLL_L_X102Y120_SLICE_X160Y120_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h90909090f00000f0)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_DLUT (
.I0(CLBLL_L_X102Y120_SLICE_X160Y120_C5Q),
.I1(CLBLL_L_X102Y121_SLICE_X161Y121_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y120_SLICE_X161Y120_B5Q),
.I4(CLBLL_L_X102Y120_SLICE_X160Y120_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y120_SLICE_X160Y120_DO5),
.O6(CLBLL_L_X102Y120_SLICE_X160Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha050a050c0c03030)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_CLUT (
.I0(CLBLL_L_X102Y119_SLICE_X160Y119_A5Q),
.I1(CLBLL_L_X102Y120_SLICE_X160Y120_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y120_SLICE_X160Y120_BQ),
.I4(CLBLL_L_X102Y119_SLICE_X160Y119_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y120_SLICE_X160Y120_CO5),
.O6(CLBLL_L_X102Y120_SLICE_X160Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00a0a28822882)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y120_SLICE_X160Y120_DQ),
.I2(CLBLM_R_X101Y117_SLICE_X159Y117_CQ),
.I3(CLBLM_R_X103Y120_SLICE_X163Y120_B5Q),
.I4(CLBLM_R_X103Y119_SLICE_X163Y119_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y120_SLICE_X160Y120_BO5),
.O6(CLBLL_L_X102Y120_SLICE_X160Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0a8888a0008888)
  ) CLBLL_L_X102Y120_SLICE_X160Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y121_SLICE_X160Y121_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X103Y120_SLICE_X162Y120_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y119_SLICE_X160Y119_DO6),
.O5(CLBLL_L_X102Y120_SLICE_X160Y120_AO5),
.O6(CLBLL_L_X102Y120_SLICE_X160Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X161Y120_BO5),
.Q(CLBLL_L_X102Y120_SLICE_X161Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X161Y120_AO6),
.Q(CLBLL_L_X102Y120_SLICE_X161Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y120_SLICE_X161Y120_BO6),
.Q(CLBLL_L_X102Y120_SLICE_X161Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699696696996)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_DLUT (
.I0(CLBLL_L_X102Y121_SLICE_X161Y121_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y120_SLICE_X161Y120_BQ),
.I3(CLBLL_L_X102Y120_SLICE_X161Y120_AQ),
.I4(CLBLL_L_X102Y120_SLICE_X161Y120_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y120_SLICE_X161Y120_DO5),
.O6(CLBLL_L_X102Y120_SLICE_X161Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a659a65959a6)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_CLUT (
.I0(CLBLL_L_X102Y121_SLICE_X161Y121_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y120_SLICE_X162Y120_A5Q),
.I3(CLBLL_L_X102Y120_SLICE_X161Y120_BQ),
.I4(CLBLL_L_X102Y120_SLICE_X161Y120_AQ),
.I5(CLBLL_L_X102Y120_SLICE_X161Y120_B5Q),
.O5(CLBLL_L_X102Y120_SLICE_X161Y120_CO5),
.O6(CLBLL_L_X102Y120_SLICE_X161Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y120_SLICE_X161Y120_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y121_SLICE_X161Y121_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y120_SLICE_X161Y120_BO5),
.O6(CLBLL_L_X102Y120_SLICE_X161Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8aaa0a8080a000)
  ) CLBLL_L_X102Y120_SLICE_X161Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y120_SLICE_X162Y120_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X102Y120_SLICE_X161Y120_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y121_SLICE_X155Y121_DO6),
.O5(CLBLL_L_X102Y120_SLICE_X161Y120_AO5),
.O6(CLBLL_L_X102Y120_SLICE_X161Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X160Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X160Y121_AO5),
.Q(CLBLL_L_X102Y121_SLICE_X160Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y121_SLICE_X160Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y121_SLICE_X160Y121_DO5),
.O6(CLBLL_L_X102Y121_SLICE_X160Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cce2e233ffe2e2)
  ) CLBLL_L_X102Y121_SLICE_X160Y121_CLUT (
.I0(CLBLM_R_X103Y125_SLICE_X162Y125_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLL_L_X102Y121_SLICE_X161Y121_DO6),
.I3(CLBLL_L_X100Y122_SLICE_X157Y122_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X102Y121_SLICE_X161Y121_C5Q),
.O5(CLBLL_L_X102Y121_SLICE_X160Y121_CO5),
.O6(CLBLL_L_X102Y121_SLICE_X160Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeeb1441ebbe4114)
  ) CLBLL_L_X102Y121_SLICE_X160Y121_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X100Y121_SLICE_X157Y121_C5Q),
.I2(CLBLL_L_X102Y121_SLICE_X160Y121_AQ),
.I3(CLBLL_L_X100Y121_SLICE_X157Y121_BQ),
.I4(CLBLL_L_X102Y120_SLICE_X160Y120_C5Q),
.I5(CLBLM_R_X101Y120_SLICE_X158Y120_CQ),
.O5(CLBLL_L_X102Y121_SLICE_X160Y121_BO5),
.O6(CLBLL_L_X102Y121_SLICE_X160Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLL_L_X102Y121_SLICE_X160Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y120_SLICE_X158Y120_CQ),
.I2(CLBLL_L_X102Y121_SLICE_X160Y121_AQ),
.I3(CLBLL_L_X100Y121_SLICE_X157Y121_BQ),
.I4(CLBLL_L_X100Y121_SLICE_X157Y121_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y121_SLICE_X160Y121_AO5),
.O6(CLBLL_L_X102Y121_SLICE_X160Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X161Y121_AO5),
.Q(CLBLL_L_X102Y121_SLICE_X161Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X161Y121_BO5),
.Q(CLBLL_L_X102Y121_SLICE_X161Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X161Y121_CO5),
.Q(CLBLL_L_X102Y121_SLICE_X161Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X161Y121_AO6),
.Q(CLBLL_L_X102Y121_SLICE_X161Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X161Y121_BO6),
.Q(CLBLL_L_X102Y121_SLICE_X161Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y121_SLICE_X161Y121_CO6),
.Q(CLBLL_L_X102Y121_SLICE_X161Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X103Y121_SLICE_X163Y121_BQ),
.I2(CLBLL_L_X102Y121_SLICE_X161Y121_BQ),
.I3(1'b1),
.I4(CLBLL_L_X102Y121_SLICE_X161Y121_B5Q),
.I5(CLBLM_R_X103Y122_SLICE_X163Y122_BQ),
.O5(CLBLL_L_X102Y121_SLICE_X161Y121_DO5),
.O6(CLBLL_L_X102Y121_SLICE_X161Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00aa00a88882222)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y121_SLICE_X161Y121_CQ),
.I2(CLBLM_R_X101Y121_SLICE_X159Y121_A5Q),
.I3(CLBLM_R_X103Y121_SLICE_X163Y121_B5Q),
.I4(CLBLL_L_X102Y121_SLICE_X161Y121_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y121_SLICE_X161Y121_CO5),
.O6(CLBLL_L_X102Y121_SLICE_X161Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y121_SLICE_X161Y121_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X103Y121_SLICE_X163Y121_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y121_SLICE_X161Y121_BO5),
.O6(CLBLL_L_X102Y121_SLICE_X161Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLL_L_X102Y121_SLICE_X161Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y120_SLICE_X161Y120_AQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y121_SLICE_X162Y121_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y121_SLICE_X161Y121_AO5),
.O6(CLBLL_L_X102Y121_SLICE_X161Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X160Y122_AO5),
.Q(CLBLL_L_X102Y122_SLICE_X160Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X160Y122_BO5),
.Q(CLBLL_L_X102Y122_SLICE_X160Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X160Y122_CO5),
.Q(CLBLL_L_X102Y122_SLICE_X160Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X160Y122_AO6),
.Q(CLBLL_L_X102Y122_SLICE_X160Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X160Y122_BO6),
.Q(CLBLL_L_X102Y122_SLICE_X160Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X160Y122_CO6),
.Q(CLBLL_L_X102Y122_SLICE_X160Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y122_SLICE_X161Y122_A5Q),
.I2(CLBLL_L_X102Y122_SLICE_X160Y122_AQ),
.I3(CLBLL_L_X102Y122_SLICE_X160Y122_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X101Y123_SLICE_X159Y123_BQ),
.O5(CLBLL_L_X102Y122_SLICE_X160Y122_DO5),
.O6(CLBLL_L_X102Y122_SLICE_X160Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0c030c030)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y122_SLICE_X161Y122_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y123_SLICE_X161Y123_A5Q),
.I4(CLBLM_R_X101Y122_SLICE_X158Y122_CO6),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X160Y122_CO5),
.O6(CLBLL_L_X102Y122_SLICE_X160Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y122_SLICE_X160Y122_B5Q),
.I2(CLBLL_L_X102Y124_SLICE_X160Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X160Y122_BO5),
.O6(CLBLL_L_X102Y122_SLICE_X160Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X102Y122_SLICE_X160Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X102Y122_SLICE_X160Y122_AQ),
.I3(CLBLM_R_X101Y123_SLICE_X159Y123_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X160Y122_AO5),
.O6(CLBLL_L_X102Y122_SLICE_X160Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X161Y122_AO5),
.Q(CLBLL_L_X102Y122_SLICE_X161Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X161Y122_BO5),
.Q(CLBLL_L_X102Y122_SLICE_X161Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X161Y122_CO5),
.Q(CLBLL_L_X102Y122_SLICE_X161Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X161Y122_AO6),
.Q(CLBLL_L_X102Y122_SLICE_X161Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X161Y122_BO6),
.Q(CLBLL_L_X102Y122_SLICE_X161Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y122_SLICE_X161Y122_CO6),
.Q(CLBLL_L_X102Y122_SLICE_X161Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X103Y123_SLICE_X162Y123_CQ),
.I2(CLBLL_L_X102Y122_SLICE_X161Y122_BQ),
.I3(CLBLL_L_X102Y122_SLICE_X161Y122_AQ),
.I4(CLBLL_L_X102Y122_SLICE_X161Y122_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X161Y122_DO5),
.O6(CLBLL_L_X102Y122_SLICE_X161Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050c0c03030)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_CLUT (
.I0(CLBLM_R_X101Y122_SLICE_X159Y122_CO6),
.I1(CLBLL_L_X102Y122_SLICE_X160Y122_C5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X102Y122_SLICE_X161Y122_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X161Y122_CO5),
.O6(CLBLL_L_X102Y122_SLICE_X161Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y122_SLICE_X161Y122_BQ),
.I2(CLBLL_L_X102Y122_SLICE_X161Y122_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X161Y122_BO5),
.O6(CLBLL_L_X102Y122_SLICE_X161Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X102Y122_SLICE_X161Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X102Y122_SLICE_X160Y122_A5Q),
.I3(CLBLM_R_X103Y123_SLICE_X162Y123_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y122_SLICE_X161Y122_AO5),
.O6(CLBLL_L_X102Y122_SLICE_X161Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y123_SLICE_X160Y123_BO5),
.Q(CLBLL_L_X102Y123_SLICE_X160Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y123_SLICE_X160Y123_AO6),
.Q(CLBLL_L_X102Y123_SLICE_X160Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y123_SLICE_X160Y123_BO6),
.Q(CLBLL_L_X102Y123_SLICE_X160Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y123_SLICE_X160Y123_AQ),
.I2(CLBLL_L_X102Y123_SLICE_X160Y123_BQ),
.I3(CLBLL_L_X102Y124_SLICE_X160Y124_CQ),
.I4(CLBLL_L_X102Y123_SLICE_X160Y123_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y123_SLICE_X160Y123_DO5),
.O6(CLBLL_L_X102Y123_SLICE_X160Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c96696996)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X102Y123_SLICE_X160Y123_AQ),
.I2(CLBLL_L_X102Y123_SLICE_X160Y123_BQ),
.I3(CLBLL_L_X102Y124_SLICE_X160Y124_CQ),
.I4(CLBLL_L_X102Y123_SLICE_X160Y123_B5Q),
.I5(CLBLL_L_X102Y122_SLICE_X160Y122_B5Q),
.O5(CLBLL_L_X102Y123_SLICE_X160Y123_CO5),
.O6(CLBLL_L_X102Y123_SLICE_X160Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y123_SLICE_X160Y123_BQ),
.I2(CLBLL_L_X102Y124_SLICE_X160Y124_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y123_SLICE_X160Y123_BO5),
.O6(CLBLL_L_X102Y123_SLICE_X160Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha808aaaaa8080000)
  ) CLBLL_L_X102Y123_SLICE_X160Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y123_SLICE_X160Y123_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y122_SLICE_X160Y122_B5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X98Y122_SLICE_X154Y122_CO6),
.O5(CLBLL_L_X102Y123_SLICE_X160Y123_AO5),
.O6(CLBLL_L_X102Y123_SLICE_X160Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y123_SLICE_X161Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y123_SLICE_X161Y123_AO5),
.Q(CLBLL_L_X102Y123_SLICE_X161Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y123_SLICE_X161Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y123_SLICE_X161Y123_AO6),
.Q(CLBLL_L_X102Y123_SLICE_X161Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h333733373f373f37)
  ) CLBLL_L_X102Y123_SLICE_X161Y123_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y122_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(1'b1),
.I5(CLBLM_R_X101Y124_SLICE_X159Y124_A5Q),
.O5(CLBLL_L_X102Y123_SLICE_X161Y123_DO5),
.O6(CLBLL_L_X102Y123_SLICE_X161Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff1dff00ff1dff)
  ) CLBLL_L_X102Y123_SLICE_X161Y123_CLUT (
.I0(RIOB33_X105Y123_IOB_X1Y123_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y123_SLICE_X161Y123_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y123_SLICE_X161Y123_CO5),
.O6(CLBLL_L_X102Y123_SLICE_X161Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h04041515ffffffff)
  ) CLBLL_L_X102Y123_SLICE_X161Y123_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y122_SLICE_X160Y122_C5Q),
.I3(1'b1),
.I4(RIOB33_X105Y123_IOB_X1Y124_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLL_L_X102Y123_SLICE_X161Y123_BO5),
.O6(CLBLL_L_X102Y123_SLICE_X161Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaa0a00a0a)
  ) CLBLL_L_X102Y123_SLICE_X161Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y124_SLICE_X159Y124_A5Q),
.I3(CLBLM_R_X101Y123_SLICE_X158Y123_CO6),
.I4(CLBLL_L_X102Y125_SLICE_X161Y125_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y123_SLICE_X161Y123_AO5),
.O6(CLBLL_L_X102Y123_SLICE_X161Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_AO5),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_CO5),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_DO5),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_AO6),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_BO6),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_CO6),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X160Y124_DO6),
.Q(CLBLL_L_X102Y124_SLICE_X160Y124_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc003300a500a500)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_DLUT (
.I0(CLBLL_L_X102Y124_SLICE_X160Y124_DQ),
.I1(CLBLL_L_X102Y124_SLICE_X161Y124_A5Q),
.I2(CLBLL_L_X102Y124_SLICE_X161Y124_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y120_SLICE_X160Y120_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y124_SLICE_X160Y124_DO5),
.O6(CLBLL_L_X102Y124_SLICE_X160Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff000000)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_CLUT (
.I0(CLBLL_L_X102Y123_SLICE_X160Y123_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X103Y124_SLICE_X163Y124_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y124_SLICE_X160Y124_CO5),
.O6(CLBLL_L_X102Y124_SLICE_X160Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88a2802200a280)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLL_L_X102Y124_SLICE_X161Y124_DO6),
.I3(CLBLM_L_X98Y123_SLICE_X154Y123_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X102Y124_SLICE_X160Y124_A5Q),
.O5(CLBLL_L_X102Y124_SLICE_X160Y124_BO5),
.O6(CLBLL_L_X102Y124_SLICE_X160Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLL_L_X102Y124_SLICE_X160Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y124_SLICE_X160Y124_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X103Y120_SLICE_X162Y120_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y124_SLICE_X160Y124_AO5),
.O6(CLBLL_L_X102Y124_SLICE_X160Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X161Y124_AO5),
.Q(CLBLL_L_X102Y124_SLICE_X161Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X161Y124_BO5),
.Q(CLBLL_L_X102Y124_SLICE_X161Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X161Y124_AO6),
.Q(CLBLL_L_X102Y124_SLICE_X161Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y124_SLICE_X161Y124_BO6),
.Q(CLBLL_L_X102Y124_SLICE_X161Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55a5aa55aa5a55a)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(1'b1),
.I2(CLBLL_L_X102Y124_SLICE_X161Y124_BQ),
.I3(CLBLL_L_X102Y124_SLICE_X161Y124_AQ),
.I4(CLBLL_L_X102Y124_SLICE_X161Y124_B5Q),
.I5(CLBLL_L_X102Y124_SLICE_X160Y124_BQ),
.O5(CLBLL_L_X102Y124_SLICE_X161Y124_DO5),
.O6(CLBLL_L_X102Y124_SLICE_X161Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22dd22d2dd2)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X102Y124_SLICE_X160Y124_A5Q),
.I2(CLBLL_L_X102Y124_SLICE_X161Y124_BQ),
.I3(CLBLL_L_X102Y124_SLICE_X161Y124_AQ),
.I4(CLBLL_L_X102Y124_SLICE_X161Y124_B5Q),
.I5(CLBLL_L_X102Y124_SLICE_X160Y124_BQ),
.O5(CLBLL_L_X102Y124_SLICE_X161Y124_CO5),
.O6(CLBLL_L_X102Y124_SLICE_X161Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y124_SLICE_X161Y124_BQ),
.I2(CLBLL_L_X102Y124_SLICE_X161Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y124_SLICE_X161Y124_BO5),
.O6(CLBLL_L_X102Y124_SLICE_X161Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X102Y124_SLICE_X161Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y124_SLICE_X162Y124_B5Q),
.I3(CLBLL_L_X102Y124_SLICE_X160Y124_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y124_SLICE_X161Y124_AO5),
.O6(CLBLL_L_X102Y124_SLICE_X161Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X160Y125_BO5),
.Q(CLBLL_L_X102Y125_SLICE_X160Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X160Y125_AO6),
.Q(CLBLL_L_X102Y125_SLICE_X160Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X160Y125_BO6),
.Q(CLBLL_L_X102Y125_SLICE_X160Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_DLUT (
.I0(CLBLM_R_X101Y126_SLICE_X159Y126_A5Q),
.I1(CLBLL_L_X102Y125_SLICE_X160Y125_AQ),
.I2(CLBLL_L_X102Y125_SLICE_X161Y125_B5Q),
.I3(CLBLL_L_X102Y125_SLICE_X160Y125_BQ),
.I4(CLBLL_L_X102Y125_SLICE_X160Y125_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_DO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_CLUT (
.I0(CLBLL_L_X102Y126_SLICE_X161Y126_AQ),
.I1(CLBLL_L_X102Y125_SLICE_X160Y125_AQ),
.I2(CLBLL_L_X102Y125_SLICE_X161Y125_B5Q),
.I3(CLBLL_L_X102Y125_SLICE_X160Y125_BQ),
.I4(CLBLL_L_X102Y125_SLICE_X160Y125_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_CO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y125_SLICE_X160Y125_BQ),
.I2(CLBLL_L_X102Y125_SLICE_X160Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_BO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa88a0000088a0)
  ) CLBLL_L_X102Y125_SLICE_X160Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_D5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y125_SLICE_X160Y125_CO6),
.O5(CLBLL_L_X102Y125_SLICE_X160Y125_AO5),
.O6(CLBLL_L_X102Y125_SLICE_X160Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X161Y125_BO5),
.Q(CLBLL_L_X102Y125_SLICE_X161Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X161Y125_CO5),
.Q(CLBLL_L_X102Y125_SLICE_X161Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X161Y125_AO6),
.Q(CLBLL_L_X102Y125_SLICE_X161Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X161Y125_BO6),
.Q(CLBLL_L_X102Y125_SLICE_X161Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y125_SLICE_X161Y125_CO6),
.Q(CLBLL_L_X102Y125_SLICE_X161Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_DLUT (
.I0(CLBLL_L_X102Y125_SLICE_X161Y125_C5Q),
.I1(CLBLL_L_X102Y125_SLICE_X161Y125_CQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y125_SLICE_X161Y125_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y125_SLICE_X161Y125_AQ),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_DO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y125_SLICE_X161Y125_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y125_SLICE_X161Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_CO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X102Y125_SLICE_X161Y125_AQ),
.I3(CLBLL_L_X102Y125_SLICE_X160Y125_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_BO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cc55ffff)
  ) CLBLL_L_X102Y125_SLICE_X161Y125_ALUT (
.I0(CLBLL_L_X102Y125_SLICE_X161Y125_DO6),
.I1(CLBLL_L_X102Y126_SLICE_X160Y126_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y123_SLICE_X161Y123_CO6),
.O5(CLBLL_L_X102Y125_SLICE_X161Y125_AO5),
.O6(CLBLL_L_X102Y125_SLICE_X161Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X160Y126_AO5),
.Q(CLBLL_L_X102Y126_SLICE_X160Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X160Y126_CO5),
.Q(CLBLL_L_X102Y126_SLICE_X160Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X160Y126_AO6),
.Q(CLBLL_L_X102Y126_SLICE_X160Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X160Y126_BO6),
.Q(CLBLL_L_X102Y126_SLICE_X160Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X160Y126_CO6),
.Q(CLBLL_L_X102Y126_SLICE_X160Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y126_SLICE_X160Y126_CQ),
.I2(CLBLL_L_X102Y126_SLICE_X160Y126_BQ),
.I3(CLBLL_L_X102Y126_SLICE_X160Y126_C5Q),
.I4(1'b1),
.I5(CLBLL_L_X102Y126_SLICE_X161Y126_C5Q),
.O5(CLBLL_L_X102Y126_SLICE_X160Y126_DO5),
.O6(CLBLL_L_X102Y126_SLICE_X160Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y126_SLICE_X160Y126_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y126_SLICE_X160Y126_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y126_SLICE_X160Y126_CO5),
.O6(CLBLL_L_X102Y126_SLICE_X160Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000f050f050f)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_BLUT (
.I0(CLBLL_L_X102Y126_SLICE_X160Y126_DO6),
.I1(1'b1),
.I2(CLBLL_L_X102Y123_SLICE_X161Y123_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLL_L_X102Y126_SLICE_X160Y126_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y126_SLICE_X160Y126_BO5),
.O6(CLBLL_L_X102Y126_SLICE_X160Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaaa0000)
  ) CLBLL_L_X102Y126_SLICE_X160Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y126_SLICE_X160Y126_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y126_SLICE_X161Y126_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y126_SLICE_X160Y126_AO5),
.O6(CLBLL_L_X102Y126_SLICE_X160Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_AO5),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_BO5),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_CO5),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_DO5),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_AO6),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_BO6),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_CO6),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y126_SLICE_X161Y126_DO6),
.Q(CLBLL_L_X102Y126_SLICE_X161Y126_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_DLUT (
.I0(CLBLL_L_X102Y126_SLICE_X161Y126_DQ),
.I1(CLBLL_L_X102Y125_SLICE_X161Y125_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X103Y126_SLICE_X162Y126_B5Q),
.I4(CLBLL_L_X102Y127_SLICE_X161Y127_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y126_SLICE_X161Y126_DO5),
.O6(CLBLL_L_X102Y126_SLICE_X161Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0c0c0c0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_CLUT (
.I0(CLBLL_L_X102Y128_SLICE_X161Y128_AQ),
.I1(CLBLL_L_X102Y126_SLICE_X160Y126_C5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y126_SLICE_X161Y126_CO5),
.O6(CLBLL_L_X102Y126_SLICE_X161Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y126_SLICE_X162Y126_AQ),
.I3(CLBLL_L_X102Y127_SLICE_X161Y127_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y126_SLICE_X161Y126_BO5),
.O6(CLBLL_L_X102Y126_SLICE_X161Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X102Y126_SLICE_X161Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_A5Q),
.I2(CLBLL_L_X102Y127_SLICE_X160Y127_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y126_SLICE_X161Y126_AO5),
.O6(CLBLL_L_X102Y126_SLICE_X161Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X160Y127_AO5),
.Q(CLBLL_L_X102Y127_SLICE_X160Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X160Y127_CO5),
.Q(CLBLL_L_X102Y127_SLICE_X160Y127_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X160Y127_AO6),
.Q(CLBLL_L_X102Y127_SLICE_X160Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X160Y127_BO6),
.Q(CLBLL_L_X102Y127_SLICE_X160Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X160Y127_CO6),
.Q(CLBLL_L_X102Y127_SLICE_X160Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006969ff009696)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_DLUT (
.I0(CLBLL_L_X102Y127_SLICE_X160Y127_C5Q),
.I1(CLBLL_L_X102Y129_SLICE_X160Y129_CQ),
.I2(CLBLL_L_X102Y127_SLICE_X160Y127_BQ),
.I3(CLBLL_L_X102Y127_SLICE_X160Y127_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X102Y127_SLICE_X160Y127_CQ),
.O5(CLBLL_L_X102Y127_SLICE_X160Y127_DO5),
.O6(CLBLL_L_X102Y127_SLICE_X160Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y127_SLICE_X160Y127_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y129_SLICE_X160Y129_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y127_SLICE_X160Y127_CO5),
.O6(CLBLL_L_X102Y127_SLICE_X160Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888aa008888a0a0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y127_SLICE_X160Y127_DO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLL_L_X102Y127_SLICE_X161Y127_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y127_SLICE_X160Y127_BO5),
.O6(CLBLL_L_X102Y127_SLICE_X160Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X102Y127_SLICE_X160Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y127_SLICE_X160Y127_A5Q),
.I2(CLBLL_L_X102Y130_SLICE_X161Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y127_SLICE_X160Y127_AO5),
.O6(CLBLL_L_X102Y127_SLICE_X160Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X161Y127_AO5),
.Q(CLBLL_L_X102Y127_SLICE_X161Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X161Y127_BO5),
.Q(CLBLL_L_X102Y127_SLICE_X161Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X161Y127_AO6),
.Q(CLBLL_L_X102Y127_SLICE_X161Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y127_SLICE_X161Y127_BO6),
.Q(CLBLL_L_X102Y127_SLICE_X161Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd8d88dd88d8dd8)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y127_SLICE_X159Y127_A5Q),
.I2(CLBLL_L_X102Y126_SLICE_X161Y126_B5Q),
.I3(CLBLL_L_X102Y127_SLICE_X161Y127_A5Q),
.I4(CLBLL_L_X102Y127_SLICE_X161Y127_AQ),
.I5(CLBLM_R_X103Y127_SLICE_X162Y127_AQ),
.O5(CLBLL_L_X102Y127_SLICE_X161Y127_DO5),
.O6(CLBLL_L_X102Y127_SLICE_X161Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_CLUT (
.I0(CLBLL_L_X102Y127_SLICE_X160Y127_AQ),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_B5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y127_SLICE_X161Y127_A5Q),
.I4(CLBLL_L_X102Y127_SLICE_X161Y127_AQ),
.I5(CLBLM_R_X103Y127_SLICE_X162Y127_AQ),
.O5(CLBLL_L_X102Y127_SLICE_X161Y127_CO5),
.O6(CLBLL_L_X102Y127_SLICE_X161Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000f0099009900)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_BLUT (
.I0(CLBLL_L_X102Y126_SLICE_X161Y126_B5Q),
.I1(CLBLL_L_X102Y127_SLICE_X161Y127_BQ),
.I2(CLBLL_L_X102Y127_SLICE_X160Y127_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y129_SLICE_X161Y129_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y127_SLICE_X161Y127_BO5),
.O6(CLBLL_L_X102Y127_SLICE_X161Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X102Y127_SLICE_X161Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X102Y127_SLICE_X161Y127_AQ),
.I3(CLBLM_R_X103Y127_SLICE_X162Y127_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y127_SLICE_X161Y127_AO5),
.O6(CLBLL_L_X102Y127_SLICE_X161Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y128_SLICE_X160Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y128_SLICE_X160Y128_DO5),
.O6(CLBLL_L_X102Y128_SLICE_X160Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y128_SLICE_X160Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y128_SLICE_X160Y128_CO5),
.O6(CLBLL_L_X102Y128_SLICE_X160Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y128_SLICE_X160Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y128_SLICE_X160Y128_BO5),
.O6(CLBLL_L_X102Y128_SLICE_X160Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y128_SLICE_X160Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y128_SLICE_X160Y128_AO5),
.O6(CLBLL_L_X102Y128_SLICE_X160Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y128_SLICE_X161Y128_BO5),
.Q(CLBLL_L_X102Y128_SLICE_X161Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y128_SLICE_X161Y128_AO6),
.Q(CLBLL_L_X102Y128_SLICE_X161Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y128_SLICE_X161Y128_BO6),
.Q(CLBLL_L_X102Y128_SLICE_X161Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_DLUT (
.I0(CLBLL_L_X102Y128_SLICE_X161Y128_BQ),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y128_SLICE_X161Y128_AQ),
.I4(CLBLL_L_X102Y128_SLICE_X161Y128_B5Q),
.I5(CLBLL_L_X100Y129_SLICE_X156Y129_AQ),
.O5(CLBLL_L_X102Y128_SLICE_X161Y128_DO5),
.O6(CLBLL_L_X102Y128_SLICE_X161Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_CLUT (
.I0(CLBLL_L_X102Y128_SLICE_X161Y128_BQ),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y128_SLICE_X161Y128_AQ),
.I4(CLBLL_L_X102Y128_SLICE_X161Y128_B5Q),
.I5(CLBLL_L_X102Y130_SLICE_X161Y130_AQ),
.O5(CLBLL_L_X102Y128_SLICE_X161Y128_CO5),
.O6(CLBLL_L_X102Y128_SLICE_X161Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y128_SLICE_X161Y128_BQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y126_SLICE_X161Y126_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y128_SLICE_X161Y128_BO5),
.O6(CLBLL_L_X102Y128_SLICE_X161Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8000000d80000)
  ) CLBLL_L_X102Y128_SLICE_X161Y128_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X102Y129_SLICE_X161Y129_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y117_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLL_L_X102Y128_SLICE_X161Y128_CO6),
.O5(CLBLL_L_X102Y128_SLICE_X161Y128_AO5),
.O6(CLBLL_L_X102Y128_SLICE_X161Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y129_SLICE_X160Y129_AO5),
.Q(CLBLL_L_X102Y129_SLICE_X160Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y129_SLICE_X160Y129_CO5),
.Q(CLBLL_L_X102Y129_SLICE_X160Y129_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y129_SLICE_X160Y129_AO6),
.Q(CLBLL_L_X102Y129_SLICE_X160Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y129_SLICE_X160Y129_BO6),
.Q(CLBLL_L_X102Y129_SLICE_X160Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y129_SLICE_X160Y129_CO6),
.Q(CLBLL_L_X102Y129_SLICE_X160Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y129_SLICE_X160Y129_DO5),
.O6(CLBLL_L_X102Y129_SLICE_X160Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ff000000)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_CLUT (
.I0(CLBLL_L_X102Y127_SLICE_X160Y127_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X102Y130_SLICE_X160Y130_B5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y129_SLICE_X160Y129_CO5),
.O6(CLBLL_L_X102Y129_SLICE_X160Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa880088aaa000a0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y130_SLICE_X161Y130_BQ),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLL_L_X102Y130_SLICE_X160Y130_CO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y129_SLICE_X160Y129_BO5),
.O6(CLBLL_L_X102Y129_SLICE_X160Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X102Y129_SLICE_X160Y129_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y129_SLICE_X160Y129_A5Q),
.I2(CLBLL_L_X100Y128_SLICE_X156Y128_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y129_SLICE_X160Y129_AO5),
.O6(CLBLL_L_X102Y129_SLICE_X160Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y129_SLICE_X161Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y129_SLICE_X161Y129_AO6),
.Q(CLBLL_L_X102Y129_SLICE_X161Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y129_SLICE_X161Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y129_SLICE_X161Y129_DO5),
.O6(CLBLL_L_X102Y129_SLICE_X161Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y129_SLICE_X161Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y129_SLICE_X161Y129_CO5),
.O6(CLBLL_L_X102Y129_SLICE_X161Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y129_SLICE_X161Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y129_SLICE_X161Y129_BO5),
.O6(CLBLL_L_X102Y129_SLICE_X161Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2288228888228822)
  ) CLBLL_L_X102Y129_SLICE_X161Y129_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y128_SLICE_X161Y128_B5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y130_SLICE_X161Y130_BQ),
.I4(1'b1),
.I5(CLBLM_R_X101Y128_SLICE_X158Y128_A5Q),
.O5(CLBLL_L_X102Y129_SLICE_X161Y129_AO5),
.O6(CLBLL_L_X102Y129_SLICE_X161Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X160Y130_AO5),
.Q(CLBLL_L_X102Y130_SLICE_X160Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X160Y130_BO5),
.Q(CLBLL_L_X102Y130_SLICE_X160Y130_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X160Y130_AO6),
.Q(CLBLL_L_X102Y130_SLICE_X160Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X160Y130_BO6),
.Q(CLBLL_L_X102Y130_SLICE_X160Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_DLUT (
.I0(CLBLL_L_X102Y129_SLICE_X160Y129_BQ),
.I1(CLBLL_L_X102Y129_SLICE_X160Y129_C5Q),
.I2(CLBLL_L_X102Y130_SLICE_X160Y130_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y130_SLICE_X160Y130_B5Q),
.I5(CLBLL_L_X100Y130_SLICE_X156Y130_AQ),
.O5(CLBLL_L_X102Y130_SLICE_X160Y130_DO5),
.O6(CLBLL_L_X102Y130_SLICE_X160Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_CLUT (
.I0(CLBLL_L_X102Y129_SLICE_X160Y129_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y129_SLICE_X160Y129_C5Q),
.I3(CLBLL_L_X102Y130_SLICE_X160Y130_BQ),
.I4(CLBLL_L_X102Y130_SLICE_X160Y130_B5Q),
.I5(CLBLL_L_X102Y130_SLICE_X161Y130_A5Q),
.O5(CLBLL_L_X102Y130_SLICE_X160Y130_CO5),
.O6(CLBLL_L_X102Y130_SLICE_X160Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y130_SLICE_X160Y130_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y129_SLICE_X160Y129_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y130_SLICE_X160Y130_BO5),
.O6(CLBLL_L_X102Y130_SLICE_X160Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888800aa00aa)
  ) CLBLL_L_X102Y130_SLICE_X160Y130_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y130_SLICE_X160Y130_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y129_SLICE_X160Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y130_SLICE_X160Y130_AO5),
.O6(CLBLL_L_X102Y130_SLICE_X160Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X161Y130_AO5),
.Q(CLBLL_L_X102Y130_SLICE_X161Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X161Y130_AO6),
.Q(CLBLL_L_X102Y130_SLICE_X161Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y130_SLICE_X161Y130_BO6),
.Q(CLBLL_L_X102Y130_SLICE_X161Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y130_SLICE_X161Y130_DO5),
.O6(CLBLL_L_X102Y130_SLICE_X161Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y130_SLICE_X161Y130_CO5),
.O6(CLBLL_L_X102Y130_SLICE_X161Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8282828282828282)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y135_SLICE_X159Y135_D5Q),
.I2(CLBLL_L_X102Y129_SLICE_X160Y129_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y130_SLICE_X161Y130_BO5),
.O6(CLBLL_L_X102Y130_SLICE_X161Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLL_L_X102Y130_SLICE_X161Y130_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y130_SLICE_X161Y130_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y134_SLICE_X160Y134_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y130_SLICE_X161Y130_AO5),
.O6(CLBLL_L_X102Y130_SLICE_X161Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y131_SLICE_X160Y131_BO5),
.Q(CLBLL_L_X102Y131_SLICE_X160Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y131_SLICE_X160Y131_AO6),
.Q(CLBLL_L_X102Y131_SLICE_X160Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y131_SLICE_X160Y131_BO6),
.Q(CLBLL_L_X102Y131_SLICE_X160Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_DLUT (
.I0(CLBLM_R_X101Y131_SLICE_X159Y131_BQ),
.I1(CLBLL_L_X102Y131_SLICE_X160Y131_AQ),
.I2(CLBLM_L_X98Y130_SLICE_X155Y130_DQ),
.I3(CLBLL_L_X102Y131_SLICE_X160Y131_BQ),
.I4(CLBLL_L_X102Y131_SLICE_X160Y131_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y131_SLICE_X160Y131_DO5),
.O6(CLBLL_L_X102Y131_SLICE_X160Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_CLUT (
.I0(CLBLM_R_X101Y131_SLICE_X159Y131_BQ),
.I1(CLBLL_L_X102Y130_SLICE_X160Y130_A5Q),
.I2(CLBLL_L_X102Y131_SLICE_X160Y131_AQ),
.I3(CLBLL_L_X102Y131_SLICE_X160Y131_BQ),
.I4(CLBLL_L_X102Y131_SLICE_X160Y131_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y131_SLICE_X160Y131_CO5),
.O6(CLBLL_L_X102Y131_SLICE_X160Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y131_SLICE_X160Y131_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y131_SLICE_X159Y131_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y131_SLICE_X160Y131_BO5),
.O6(CLBLL_L_X102Y131_SLICE_X160Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa2a8a00a020800)
  ) CLBLL_L_X102Y131_SLICE_X160Y131_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y131_SLICE_X159Y131_CQ),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLL_L_X102Y131_SLICE_X160Y131_CO6),
.O5(CLBLL_L_X102Y131_SLICE_X160Y131_AO5),
.O6(CLBLL_L_X102Y131_SLICE_X160Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y131_SLICE_X161Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y131_SLICE_X161Y131_DO5),
.O6(CLBLL_L_X102Y131_SLICE_X161Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y131_SLICE_X161Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y131_SLICE_X161Y131_CO5),
.O6(CLBLL_L_X102Y131_SLICE_X161Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y131_SLICE_X161Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y131_SLICE_X161Y131_BO5),
.O6(CLBLL_L_X102Y131_SLICE_X161Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y131_SLICE_X161Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y131_SLICE_X161Y131_AO5),
.O6(CLBLL_L_X102Y131_SLICE_X161Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y134_SLICE_X160Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y134_SLICE_X160Y134_AO5),
.Q(CLBLL_L_X102Y134_SLICE_X160Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y134_SLICE_X160Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y134_SLICE_X160Y134_AO6),
.Q(CLBLL_L_X102Y134_SLICE_X160Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X160Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X160Y134_DO5),
.O6(CLBLL_L_X102Y134_SLICE_X160Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X160Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X160Y134_CO5),
.O6(CLBLL_L_X102Y134_SLICE_X160Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X160Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X160Y134_BO5),
.O6(CLBLL_L_X102Y134_SLICE_X160Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLL_L_X102Y134_SLICE_X160Y134_ALUT (
.I0(CLBLM_R_X101Y136_SLICE_X158Y136_AQ),
.I1(CLBLL_L_X102Y134_SLICE_X160Y134_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X160Y134_AO5),
.O6(CLBLL_L_X102Y134_SLICE_X160Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X161Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X161Y134_DO5),
.O6(CLBLL_L_X102Y134_SLICE_X161Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X161Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X161Y134_CO5),
.O6(CLBLL_L_X102Y134_SLICE_X161Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X161Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X161Y134_BO5),
.O6(CLBLL_L_X102Y134_SLICE_X161Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y134_SLICE_X161Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y134_SLICE_X161Y134_AO5),
.O6(CLBLL_L_X102Y134_SLICE_X161Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y135_SLICE_X160Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y135_SLICE_X160Y135_AO6),
.Q(CLBLL_L_X102Y135_SLICE_X160Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y135_SLICE_X160Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y135_SLICE_X160Y135_DO5),
.O6(CLBLL_L_X102Y135_SLICE_X160Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLL_L_X102Y135_SLICE_X160Y135_CLUT (
.I0(CLBLL_L_X102Y136_SLICE_X160Y136_AQ),
.I1(CLBLL_L_X100Y134_SLICE_X156Y134_B5Q),
.I2(CLBLL_L_X102Y136_SLICE_X160Y136_BQ),
.I3(CLBLM_R_X101Y135_SLICE_X159Y135_BQ),
.I4(CLBLL_L_X102Y136_SLICE_X160Y136_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLL_L_X102Y135_SLICE_X160Y135_CO5),
.O6(CLBLL_L_X102Y135_SLICE_X160Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLL_L_X102Y135_SLICE_X160Y135_BLUT (
.I0(CLBLM_R_X101Y135_SLICE_X158Y135_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y135_SLICE_X160Y135_AQ),
.I3(CLBLM_R_X101Y135_SLICE_X159Y135_AQ),
.I4(CLBLL_L_X102Y134_SLICE_X160Y134_AQ),
.I5(CLBLM_R_X101Y135_SLICE_X158Y135_AQ),
.O5(CLBLL_L_X102Y135_SLICE_X160Y135_BO5),
.O6(CLBLL_L_X102Y135_SLICE_X160Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa5000000000)
  ) CLBLL_L_X102Y135_SLICE_X160Y135_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y135_SLICE_X159Y135_D5Q),
.I2(RIOB33_X105Y145_IOB_X1Y145_I),
.I3(CLBLL_L_X102Y135_SLICE_X160Y135_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLL_L_X102Y135_SLICE_X160Y135_AO5),
.O6(CLBLL_L_X102Y135_SLICE_X160Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y135_SLICE_X161Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y135_SLICE_X161Y135_DO5),
.O6(CLBLL_L_X102Y135_SLICE_X161Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y135_SLICE_X161Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y135_SLICE_X161Y135_CO5),
.O6(CLBLL_L_X102Y135_SLICE_X161Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y135_SLICE_X161Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y135_SLICE_X161Y135_BO5),
.O6(CLBLL_L_X102Y135_SLICE_X161Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y135_SLICE_X161Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y135_SLICE_X161Y135_AO5),
.O6(CLBLL_L_X102Y135_SLICE_X161Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y136_SLICE_X160Y136_BO5),
.Q(CLBLL_L_X102Y136_SLICE_X160Y136_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y136_SLICE_X160Y136_AO6),
.Q(CLBLL_L_X102Y136_SLICE_X160Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y136_SLICE_X160Y136_BO6),
.Q(CLBLL_L_X102Y136_SLICE_X160Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y136_SLICE_X160Y136_DO5),
.O6(CLBLL_L_X102Y136_SLICE_X160Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_CLUT (
.I0(CLBLL_L_X102Y136_SLICE_X160Y136_BQ),
.I1(CLBLL_L_X102Y136_SLICE_X160Y136_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X101Y135_SLICE_X159Y135_BQ),
.I4(CLBLL_L_X102Y136_SLICE_X160Y136_B5Q),
.I5(CLBLM_R_X101Y136_SLICE_X158Y136_AQ),
.O5(CLBLL_L_X102Y136_SLICE_X160Y136_CO5),
.O6(CLBLL_L_X102Y136_SLICE_X160Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_BLUT (
.I0(CLBLM_R_X101Y135_SLICE_X159Y135_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y136_SLICE_X160Y136_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y136_SLICE_X160Y136_BO5),
.O6(CLBLL_L_X102Y136_SLICE_X160Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e0200000e020)
  ) CLBLL_L_X102Y136_SLICE_X160Y136_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y135_SLICE_X159Y135_C5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X102Y136_SLICE_X160Y136_CO6),
.O5(CLBLL_L_X102Y136_SLICE_X160Y136_AO5),
.O6(CLBLL_L_X102Y136_SLICE_X160Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y136_SLICE_X161Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y136_SLICE_X161Y136_DO5),
.O6(CLBLL_L_X102Y136_SLICE_X161Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y136_SLICE_X161Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y136_SLICE_X161Y136_CO5),
.O6(CLBLL_L_X102Y136_SLICE_X161Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y136_SLICE_X161Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y136_SLICE_X161Y136_BO5),
.O6(CLBLL_L_X102Y136_SLICE_X161Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y136_SLICE_X161Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y136_SLICE_X161Y136_AO5),
.O6(CLBLL_L_X102Y136_SLICE_X161Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_R_X87Y118_SLICE_X138Y118_BO5),
.Q(CLBLL_R_X87Y118_SLICE_X138Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_R_X87Y118_SLICE_X138Y118_AO5),
.Q(CLBLL_R_X87Y118_SLICE_X138Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_R_X87Y118_SLICE_X138Y118_BO6),
.Q(CLBLL_R_X87Y118_SLICE_X138Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X87Y118_SLICE_X138Y118_DO5),
.O6(CLBLL_R_X87Y118_SLICE_X138Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X87Y118_SLICE_X138Y118_CO5),
.O6(CLBLL_R_X87Y118_SLICE_X138Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_BLUT (
.I0(1'b1),
.I1(CLBLL_R_X87Y118_SLICE_X138Y118_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_R_X87Y118_SLICE_X139Y118_AQ),
.I5(1'b1),
.O5(CLBLL_R_X87Y118_SLICE_X138Y118_BO5),
.O6(CLBLL_R_X87Y118_SLICE_X138Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caa00aa00)
  ) CLBLL_R_X87Y118_SLICE_X138Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_R_X87Y118_SLICE_X138Y118_BQ),
.I2(CLBLL_R_X87Y118_SLICE_X138Y118_AQ),
.I3(CLBLL_R_X87Y118_SLICE_X138Y118_B5Q),
.I4(CLBLL_R_X87Y118_SLICE_X139Y118_AQ),
.I5(1'b1),
.O5(CLBLL_R_X87Y118_SLICE_X138Y118_AO5),
.O6(CLBLL_R_X87Y118_SLICE_X138Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X87Y118_SLICE_X139Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_R_X87Y118_SLICE_X139Y118_AO6),
.Q(CLBLL_R_X87Y118_SLICE_X139Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X87Y118_SLICE_X139Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X87Y118_SLICE_X139Y118_DO5),
.O6(CLBLL_R_X87Y118_SLICE_X139Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X87Y118_SLICE_X139Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X87Y118_SLICE_X139Y118_CO5),
.O6(CLBLL_R_X87Y118_SLICE_X139Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd8d88dd88d8dd8)
  ) CLBLL_R_X87Y118_SLICE_X139Y118_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X89Y118_SLICE_X141Y118_DQ),
.I2(CLBLL_R_X87Y118_SLICE_X139Y118_AQ),
.I3(CLBLL_R_X87Y118_SLICE_X138Y118_BQ),
.I4(CLBLL_R_X87Y118_SLICE_X138Y118_AQ),
.I5(CLBLL_R_X87Y118_SLICE_X138Y118_B5Q),
.O5(CLBLL_R_X87Y118_SLICE_X139Y118_BO5),
.O6(CLBLL_R_X87Y118_SLICE_X139Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaa30aa00000000)
  ) CLBLL_R_X87Y118_SLICE_X139Y118_ALUT (
.I0(CLBLM_R_X89Y121_SLICE_X141Y121_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_R_X87Y118_SLICE_X138Y118_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X89Y119_SLICE_X140Y119_BQ),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLL_R_X87Y118_SLICE_X139Y118_AO5),
.O6(CLBLL_R_X87Y118_SLICE_X139Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X142Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X142Y113_AO5),
.Q(CLBLM_L_X90Y113_SLICE_X142Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X142Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X142Y113_AO6),
.Q(CLBLM_L_X90Y113_SLICE_X142Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y113_SLICE_X142Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y113_SLICE_X142Y113_DO5),
.O6(CLBLM_L_X90Y113_SLICE_X142Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X90Y113_SLICE_X142Y113_CLUT (
.I0(CLBLM_L_X90Y113_SLICE_X143Y113_AQ),
.I1(1'b1),
.I2(CLBLM_L_X90Y113_SLICE_X142Y113_AQ),
.I3(CLBLM_L_X90Y113_SLICE_X142Y113_A5Q),
.I4(CLBLM_L_X90Y114_SLICE_X143Y114_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X90Y113_SLICE_X142Y113_CO5),
.O6(CLBLM_L_X90Y113_SLICE_X142Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h54f45efe04a40eae)
  ) CLBLM_L_X90Y113_SLICE_X142Y113_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X92Y114_SLICE_X144Y114_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X90Y114_SLICE_X142Y114_B5Q),
.I4(CLBLM_L_X92Y115_SLICE_X145Y115_B5Q),
.I5(CLBLM_L_X90Y113_SLICE_X142Y113_CO6),
.O5(CLBLM_L_X90Y113_SLICE_X142Y113_BO5),
.O6(CLBLM_L_X90Y113_SLICE_X142Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_L_X90Y113_SLICE_X142Y113_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X90Y113_SLICE_X142Y113_AQ),
.I3(1'b1),
.I4(CLBLM_L_X90Y113_SLICE_X143Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y113_SLICE_X142Y113_AO5),
.O6(CLBLM_L_X90Y113_SLICE_X142Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X143Y113_AO5),
.Q(CLBLM_L_X90Y113_SLICE_X143Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X143Y113_BO5),
.Q(CLBLM_L_X90Y113_SLICE_X143Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X143Y113_CO5),
.Q(CLBLM_L_X90Y113_SLICE_X143Y113_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X143Y113_AO6),
.Q(CLBLM_L_X90Y113_SLICE_X143Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X143Y113_BO6),
.Q(CLBLM_L_X90Y113_SLICE_X143Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y113_SLICE_X143Y113_CO6),
.Q(CLBLM_L_X90Y113_SLICE_X143Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_DLUT (
.I0(CLBLM_L_X90Y113_SLICE_X143Y113_C5Q),
.I1(CLBLM_L_X90Y113_SLICE_X143Y113_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X90Y113_SLICE_X143Y113_B5Q),
.I5(CLBLM_R_X93Y114_SLICE_X146Y114_BQ),
.O5(CLBLM_L_X90Y113_SLICE_X143Y113_DO5),
.O6(CLBLM_L_X90Y113_SLICE_X143Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y113_SLICE_X143Y113_CQ),
.I2(1'b1),
.I3(CLBLM_R_X93Y114_SLICE_X146Y114_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y113_SLICE_X143Y113_CO5),
.O6(CLBLM_L_X90Y113_SLICE_X143Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y114_SLICE_X146Y114_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y113_SLICE_X143Y113_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y113_SLICE_X143Y113_BO5),
.O6(CLBLM_L_X90Y113_SLICE_X143Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300aa005500)
  ) CLBLM_L_X90Y113_SLICE_X143Y113_ALUT (
.I0(CLBLM_L_X90Y113_SLICE_X143Y113_B5Q),
.I1(CLBLM_L_X90Y113_SLICE_X142Y113_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y113_SLICE_X145Y113_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y113_SLICE_X143Y113_AO5),
.O6(CLBLM_L_X90Y113_SLICE_X143Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X142Y114_AO5),
.Q(CLBLM_L_X90Y114_SLICE_X142Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X142Y114_BO5),
.Q(CLBLM_L_X90Y114_SLICE_X142Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X142Y114_CO5),
.Q(CLBLM_L_X90Y114_SLICE_X142Y114_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X142Y114_AO6),
.Q(CLBLM_L_X90Y114_SLICE_X142Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X142Y114_BO6),
.Q(CLBLM_L_X90Y114_SLICE_X142Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X142Y114_CO6),
.Q(CLBLM_L_X90Y114_SLICE_X142Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_DLUT (
.I0(CLBLM_L_X90Y114_SLICE_X142Y114_C5Q),
.I1(CLBLM_L_X90Y114_SLICE_X142Y114_CQ),
.I2(CLBLM_R_X89Y114_SLICE_X141Y114_A5Q),
.I3(CLBLM_L_X90Y115_SLICE_X143Y115_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y114_SLICE_X142Y114_DO5),
.O6(CLBLM_L_X90Y114_SLICE_X142Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y114_SLICE_X142Y114_CQ),
.I2(1'b1),
.I3(CLBLM_L_X90Y115_SLICE_X143Y115_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y114_SLICE_X142Y114_CO5),
.O6(CLBLM_L_X90Y114_SLICE_X142Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000cccc0000)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_BLUT (
.I0(CLBLM_L_X90Y114_SLICE_X142Y114_B5Q),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y114_SLICE_X142Y114_BO5),
.O6(CLBLM_L_X90Y114_SLICE_X142Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00000f0f0000)
  ) CLBLM_L_X90Y114_SLICE_X142Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y114_SLICE_X142Y114_BQ),
.I2(CLBLM_L_X90Y114_SLICE_X142Y114_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y114_SLICE_X142Y114_AO5),
.O6(CLBLM_L_X90Y114_SLICE_X142Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X143Y114_AO5),
.Q(CLBLM_L_X90Y114_SLICE_X143Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X143Y114_BO5),
.Q(CLBLM_L_X90Y114_SLICE_X143Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X143Y114_AO6),
.Q(CLBLM_L_X90Y114_SLICE_X143Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y114_SLICE_X143Y114_BO6),
.Q(CLBLM_L_X90Y114_SLICE_X143Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_DLUT (
.I0(CLBLM_L_X90Y114_SLICE_X143Y114_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X90Y114_SLICE_X143Y114_AQ),
.I4(CLBLM_L_X90Y114_SLICE_X143Y114_B5Q),
.I5(CLBLM_L_X92Y114_SLICE_X144Y114_AQ),
.O5(CLBLM_L_X90Y114_SLICE_X143Y114_DO5),
.O6(CLBLM_L_X90Y114_SLICE_X143Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h323e020ef2fec2ce)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_CLUT (
.I0(CLBLM_L_X90Y118_SLICE_X143Y118_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X90Y115_SLICE_X143Y115_B5Q),
.I4(CLBLM_L_X90Y114_SLICE_X143Y114_DO6),
.I5(CLBLM_L_X90Y114_SLICE_X142Y114_BQ),
.O5(CLBLM_L_X90Y114_SLICE_X143Y114_CO5),
.O6(CLBLM_L_X90Y114_SLICE_X143Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0c0c0c0)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_BLUT (
.I0(CLBLM_L_X90Y114_SLICE_X143Y114_AQ),
.I1(CLBLM_L_X90Y114_SLICE_X143Y114_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y114_SLICE_X143Y114_BO5),
.O6(CLBLM_L_X90Y114_SLICE_X143Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000a0a0a0a0)
  ) CLBLM_L_X90Y114_SLICE_X143Y114_ALUT (
.I0(CLBLM_L_X90Y113_SLICE_X142Y113_A5Q),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X92Y114_SLICE_X144Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y114_SLICE_X143Y114_AO5),
.O6(CLBLM_L_X90Y114_SLICE_X143Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X142Y115_AO5),
.Q(CLBLM_L_X90Y115_SLICE_X142Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X142Y115_AO6),
.Q(CLBLM_L_X90Y115_SLICE_X142Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X142Y115_BO6),
.Q(CLBLM_L_X90Y115_SLICE_X142Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y115_SLICE_X142Y115_DO5),
.O6(CLBLM_L_X90Y115_SLICE_X142Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3175b9fd2064a8ec)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X90Y114_SLICE_X142Y114_DO6),
.I3(CLBLM_L_X90Y115_SLICE_X142Y115_A5Q),
.I4(CLBLM_L_X90Y114_SLICE_X142Y114_AQ),
.I5(CLBLM_L_X90Y117_SLICE_X143Y117_DO6),
.O5(CLBLM_L_X90Y115_SLICE_X142Y115_CO5),
.O6(CLBLM_L_X90Y115_SLICE_X142Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he040f0f0e0400000)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X90Y116_SLICE_X142Y116_BO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y117_SLICE_X140Y117_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X89Y115_SLICE_X140Y115_DO6),
.O5(CLBLM_L_X90Y115_SLICE_X142Y115_BO5),
.O6(CLBLM_L_X90Y115_SLICE_X142Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030a0a05050)
  ) CLBLM_L_X90Y115_SLICE_X142Y115_ALUT (
.I0(CLBLM_L_X90Y115_SLICE_X143Y115_B5Q),
.I1(CLBLM_L_X90Y115_SLICE_X143Y115_DO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X89Y114_SLICE_X141Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y115_SLICE_X142Y115_AO5),
.O6(CLBLM_L_X90Y115_SLICE_X142Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X143Y115_AO5),
.Q(CLBLM_L_X90Y115_SLICE_X143Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X143Y115_BO5),
.Q(CLBLM_L_X90Y115_SLICE_X143Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X143Y115_CO5),
.Q(CLBLM_L_X90Y115_SLICE_X143Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X143Y115_AO6),
.Q(CLBLM_L_X90Y115_SLICE_X143Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X143Y115_BO6),
.Q(CLBLM_L_X90Y115_SLICE_X143Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y115_SLICE_X143Y115_CO6),
.Q(CLBLM_L_X90Y115_SLICE_X143Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0afa0c0c0afafcfc)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_DLUT (
.I0(CLBLM_R_X89Y115_SLICE_X141Y115_DO6),
.I1(CLBLM_R_X89Y114_SLICE_X141Y114_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y115_SLICE_X143Y115_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X89Y115_SLICE_X141Y115_CQ),
.O5(CLBLM_L_X90Y115_SLICE_X143Y115_DO5),
.O6(CLBLM_L_X90Y115_SLICE_X143Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y115_SLICE_X142Y115_CO6),
.I2(CLBLM_L_X92Y114_SLICE_X144Y114_A5Q),
.I3(CLBLM_L_X90Y117_SLICE_X143Y117_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y115_SLICE_X143Y115_CO5),
.O6(CLBLM_L_X90Y115_SLICE_X143Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050c030c030)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_BLUT (
.I0(CLBLM_L_X92Y115_SLICE_X145Y115_CO6),
.I1(CLBLM_L_X90Y114_SLICE_X143Y114_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y115_SLICE_X145Y115_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y115_SLICE_X143Y115_BO5),
.O6(CLBLM_L_X90Y115_SLICE_X143Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X90Y115_SLICE_X143Y115_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y117_SLICE_X140Y117_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y115_SLICE_X143Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y115_SLICE_X143Y115_AO5),
.O6(CLBLM_L_X90Y115_SLICE_X143Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X142Y116_AO5),
.Q(CLBLM_L_X90Y116_SLICE_X142Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X142Y116_CO5),
.Q(CLBLM_L_X90Y116_SLICE_X142Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X142Y116_AO6),
.Q(CLBLM_L_X90Y116_SLICE_X142Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X142Y116_BO5),
.Q(CLBLM_L_X90Y116_SLICE_X142Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X142Y116_CO6),
.Q(CLBLM_L_X90Y116_SLICE_X142Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cacac5cac5c5ca)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_DLUT (
.I0(CLBLM_L_X90Y116_SLICE_X142Y116_C5Q),
.I1(CLBLM_R_X95Y117_SLICE_X150Y117_C5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y116_SLICE_X142Y116_BQ),
.I4(CLBLM_L_X90Y117_SLICE_X142Y117_CQ),
.I5(CLBLM_L_X90Y115_SLICE_X142Y115_BQ),
.O5(CLBLM_L_X90Y116_SLICE_X142Y116_DO5),
.O6(CLBLM_L_X90Y116_SLICE_X142Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X90Y116_SLICE_X142Y116_AQ),
.I3(1'b1),
.I4(CLBLM_L_X90Y117_SLICE_X142Y117_CQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y116_SLICE_X142Y116_CO5),
.O6(CLBLM_L_X90Y116_SLICE_X142Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_BLUT (
.I0(CLBLM_L_X90Y117_SLICE_X142Y117_CQ),
.I1(CLBLM_L_X90Y116_SLICE_X142Y116_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y115_SLICE_X142Y115_BQ),
.I4(CLBLM_L_X90Y116_SLICE_X142Y116_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y116_SLICE_X142Y116_BO5),
.O6(CLBLM_L_X90Y116_SLICE_X142Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000066990000)
  ) CLBLM_L_X90Y116_SLICE_X142Y116_ALUT (
.I0(CLBLM_R_X89Y114_SLICE_X141Y114_B5Q),
.I1(CLBLM_L_X90Y115_SLICE_X142Y115_A5Q),
.I2(CLBLM_L_X92Y116_SLICE_X145Y116_CO6),
.I3(CLBLM_L_X90Y119_SLICE_X142Y119_C5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y116_SLICE_X142Y116_AO5),
.O6(CLBLM_L_X90Y116_SLICE_X142Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X143Y116_AO5),
.Q(CLBLM_L_X90Y116_SLICE_X143Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X143Y116_BO5),
.Q(CLBLM_L_X90Y116_SLICE_X143Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X143Y116_CO5),
.Q(CLBLM_L_X90Y116_SLICE_X143Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X143Y116_AO6),
.Q(CLBLM_L_X90Y116_SLICE_X143Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X143Y116_BO6),
.Q(CLBLM_L_X90Y116_SLICE_X143Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y116_SLICE_X143Y116_CO6),
.Q(CLBLM_L_X90Y116_SLICE_X143Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303fa0af3f3fa0a)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_DLUT (
.I0(CLBLM_L_X92Y120_SLICE_X144Y120_DO6),
.I1(CLBLM_L_X90Y116_SLICE_X142Y116_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X89Y114_SLICE_X141Y114_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y116_SLICE_X140Y116_AQ),
.O5(CLBLM_L_X90Y116_SLICE_X143Y116_DO5),
.O6(CLBLM_L_X90Y116_SLICE_X143Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88228822a0a00a0a)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y116_SLICE_X142Y116_A5Q),
.I2(CLBLM_L_X92Y116_SLICE_X144Y116_B5Q),
.I3(CLBLM_L_X92Y116_SLICE_X144Y116_A5Q),
.I4(CLBLM_L_X90Y116_SLICE_X143Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y116_SLICE_X143Y116_CO5),
.O6(CLBLM_L_X90Y116_SLICE_X143Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050c030c030)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_BLUT (
.I0(CLBLM_L_X90Y116_SLICE_X143Y116_DO6),
.I1(CLBLM_L_X90Y115_SLICE_X143Y115_C5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y117_SLICE_X143Y117_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y116_SLICE_X143Y116_BO5),
.O6(CLBLM_L_X90Y116_SLICE_X143Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X90Y116_SLICE_X143Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y116_SLICE_X140Y116_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y116_SLICE_X143Y116_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y116_SLICE_X143Y116_AO5),
.O6(CLBLM_L_X90Y116_SLICE_X143Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X142Y117_BO5),
.Q(CLBLM_L_X90Y117_SLICE_X142Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X142Y117_CO5),
.Q(CLBLM_L_X90Y117_SLICE_X142Y117_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X142Y117_AO6),
.Q(CLBLM_L_X90Y117_SLICE_X142Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X142Y117_CO6),
.Q(CLBLM_L_X90Y117_SLICE_X142Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_DLUT (
.I0(CLBLM_L_X90Y117_SLICE_X142Y117_C5Q),
.I1(CLBLM_L_X90Y117_SLICE_X142Y117_AQ),
.I2(CLBLM_R_X95Y117_SLICE_X150Y117_CQ),
.I3(CLBLM_L_X90Y117_SLICE_X142Y117_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X90Y119_SLICE_X142Y119_BQ),
.O5(CLBLM_L_X90Y117_SLICE_X142Y117_DO5),
.O6(CLBLM_L_X90Y117_SLICE_X142Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X90Y119_SLICE_X142Y119_BQ),
.I3(1'b1),
.I4(CLBLM_L_X90Y115_SLICE_X142Y115_BQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y117_SLICE_X142Y117_CO5),
.O6(CLBLM_L_X90Y117_SLICE_X142Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_BLUT (
.I0(CLBLM_L_X90Y117_SLICE_X142Y117_AQ),
.I1(CLBLM_L_X90Y117_SLICE_X142Y117_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y119_SLICE_X142Y119_BQ),
.I4(CLBLM_L_X90Y117_SLICE_X142Y117_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y117_SLICE_X142Y117_BO5),
.O6(CLBLM_L_X90Y117_SLICE_X142Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d80000fa500000)
  ) CLBLM_L_X90Y117_SLICE_X142Y117_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X89Y117_SLICE_X140Y117_A5Q),
.I2(CLBLM_R_X89Y116_SLICE_X141Y116_DO6),
.I3(CLBLM_L_X90Y117_SLICE_X142Y117_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y117_SLICE_X142Y117_AO5),
.O6(CLBLM_L_X90Y117_SLICE_X142Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X143Y117_AO5),
.Q(CLBLM_L_X90Y117_SLICE_X143Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X143Y117_BO5),
.Q(CLBLM_L_X90Y117_SLICE_X143Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X143Y117_AO6),
.Q(CLBLM_L_X90Y117_SLICE_X143Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y117_SLICE_X143Y117_BO6),
.Q(CLBLM_L_X90Y117_SLICE_X143Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_DLUT (
.I0(CLBLM_L_X90Y117_SLICE_X143Y117_BQ),
.I1(CLBLM_L_X90Y117_SLICE_X143Y117_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y119_SLICE_X146Y119_AQ),
.I4(CLBLM_L_X90Y117_SLICE_X143Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y117_SLICE_X143Y117_DO5),
.O6(CLBLM_L_X90Y117_SLICE_X143Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h777730fc444430fc)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_CLUT (
.I0(CLBLM_L_X90Y116_SLICE_X143Y116_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X92Y119_SLICE_X145Y119_DO6),
.I3(CLBLM_L_X90Y116_SLICE_X143Y116_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X90Y118_SLICE_X142Y118_DO6),
.O5(CLBLM_L_X90Y117_SLICE_X143Y117_CO5),
.O6(CLBLM_L_X90Y117_SLICE_X143Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y117_SLICE_X143Y117_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y117_SLICE_X143Y117_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y117_SLICE_X143Y117_BO5),
.O6(CLBLM_L_X90Y117_SLICE_X143Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f0f00000)
  ) CLBLM_L_X90Y117_SLICE_X143Y117_ALUT (
.I0(CLBLM_R_X93Y119_SLICE_X146Y119_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y118_SLICE_X143Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y117_SLICE_X143Y117_AO5),
.O6(CLBLM_L_X90Y117_SLICE_X143Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X142Y118_AO5),
.Q(CLBLM_L_X90Y118_SLICE_X142Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X142Y118_BO5),
.Q(CLBLM_L_X90Y118_SLICE_X142Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X142Y118_AO6),
.Q(CLBLM_L_X90Y118_SLICE_X142Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X142Y118_BO6),
.Q(CLBLM_L_X90Y118_SLICE_X142Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_DLUT (
.I0(CLBLM_L_X90Y120_SLICE_X143Y120_AQ),
.I1(CLBLM_L_X92Y116_SLICE_X144Y116_A5Q),
.I2(CLBLM_L_X90Y118_SLICE_X142Y118_BQ),
.I3(1'b1),
.I4(CLBLM_L_X90Y118_SLICE_X142Y118_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X90Y118_SLICE_X142Y118_DO5),
.O6(CLBLM_L_X90Y118_SLICE_X142Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3cc3aaaac33c)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_CLUT (
.I0(CLBLM_R_X95Y118_SLICE_X150Y118_CQ),
.I1(CLBLM_R_X89Y118_SLICE_X140Y118_BQ),
.I2(CLBLM_R_X89Y118_SLICE_X140Y118_B5Q),
.I3(CLBLM_L_X90Y118_SLICE_X142Y118_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y118_SLICE_X140Y118_DQ),
.O5(CLBLM_L_X90Y118_SLICE_X142Y118_CO5),
.O6(CLBLM_L_X90Y118_SLICE_X142Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y118_SLICE_X142Y118_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y120_SLICE_X143Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y118_SLICE_X142Y118_BO5),
.O6(CLBLM_L_X90Y118_SLICE_X142Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0a0a0a0a0)
  ) CLBLM_L_X90Y118_SLICE_X142Y118_ALUT (
.I0(CLBLM_R_X89Y118_SLICE_X140Y118_DQ),
.I1(CLBLM_R_X89Y117_SLICE_X140Y117_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y118_SLICE_X142Y118_AO5),
.O6(CLBLM_L_X90Y118_SLICE_X142Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X143Y118_AO5),
.Q(CLBLM_L_X90Y118_SLICE_X143Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X143Y118_BO5),
.Q(CLBLM_L_X90Y118_SLICE_X143Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X143Y118_AO6),
.Q(CLBLM_L_X90Y118_SLICE_X143Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y118_SLICE_X143Y118_BO6),
.Q(CLBLM_L_X90Y118_SLICE_X143Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X90Y117_SLICE_X143Y117_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X90Y118_SLICE_X143Y118_BQ),
.I4(CLBLM_L_X90Y118_SLICE_X143Y118_B5Q),
.I5(CLBLM_R_X93Y119_SLICE_X146Y119_BQ),
.O5(CLBLM_L_X90Y118_SLICE_X143Y118_DO5),
.O6(CLBLM_L_X90Y118_SLICE_X143Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11ddfcfc11dd3030)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_CLUT (
.I0(CLBLM_L_X90Y115_SLICE_X143Y115_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X93Y119_SLICE_X146Y119_DO6),
.I3(CLBLM_L_X90Y118_SLICE_X143Y118_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X90Y118_SLICE_X143Y118_DO6),
.O5(CLBLM_L_X90Y118_SLICE_X143Y118_CO5),
.O6(CLBLM_L_X90Y118_SLICE_X143Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y118_SLICE_X143Y118_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y119_SLICE_X146Y119_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y118_SLICE_X143Y118_BO5),
.O6(CLBLM_L_X90Y118_SLICE_X143Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0a0a0a0a0)
  ) CLBLM_L_X90Y118_SLICE_X143Y118_ALUT (
.I0(CLBLM_L_X92Y114_SLICE_X145Y114_AQ),
.I1(CLBLM_L_X90Y118_SLICE_X143Y118_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y118_SLICE_X143Y118_AO5),
.O6(CLBLM_L_X90Y118_SLICE_X143Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X142Y119_BO5),
.Q(CLBLM_L_X90Y119_SLICE_X142Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X142Y119_CO5),
.Q(CLBLM_L_X90Y119_SLICE_X142Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X142Y119_BO6),
.Q(CLBLM_L_X90Y119_SLICE_X142Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X142Y119_CO6),
.Q(CLBLM_L_X90Y119_SLICE_X142Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5acca5cca5cc5a)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_DLUT (
.I0(CLBLM_L_X90Y119_SLICE_X143Y119_AQ),
.I1(CLBLM_R_X95Y118_SLICE_X150Y118_C5Q),
.I2(CLBLM_L_X90Y118_SLICE_X142Y118_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X90Y119_SLICE_X142Y119_B5Q),
.I5(CLBLM_R_X89Y117_SLICE_X140Y117_BQ),
.O5(CLBLM_L_X90Y119_SLICE_X142Y119_DO5),
.O6(CLBLM_L_X90Y119_SLICE_X142Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88228822a0a00a0a)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y120_SLICE_X141Y120_C5Q),
.I2(CLBLM_R_X89Y115_SLICE_X140Y115_A5Q),
.I3(CLBLM_R_X89Y116_SLICE_X140Y116_B5Q),
.I4(CLBLM_L_X90Y119_SLICE_X142Y119_CQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y119_SLICE_X142Y119_CO5),
.O6(CLBLM_L_X90Y119_SLICE_X142Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y118_SLICE_X142Y118_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y117_SLICE_X142Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y119_SLICE_X142Y119_BO5),
.O6(CLBLM_L_X90Y119_SLICE_X142Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_L_X90Y119_SLICE_X142Y119_ALUT (
.I0(CLBLM_L_X90Y119_SLICE_X142Y119_B5Q),
.I1(CLBLM_R_X89Y117_SLICE_X140Y117_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y118_SLICE_X142Y118_AQ),
.I4(CLBLM_L_X90Y119_SLICE_X143Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y119_SLICE_X142Y119_AO5),
.O6(CLBLM_L_X90Y119_SLICE_X142Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X143Y119_BO5),
.Q(CLBLM_L_X90Y119_SLICE_X143Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X142Y119_AO5),
.Q(CLBLM_L_X90Y119_SLICE_X143Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X143Y119_BO6),
.Q(CLBLM_L_X90Y119_SLICE_X143Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y119_SLICE_X143Y119_AO5),
.Q(CLBLM_L_X90Y119_SLICE_X143Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1b1b1b1bffaa5500)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X90Y116_SLICE_X143Y116_B5Q),
.I2(CLBLM_L_X90Y118_SLICE_X143Y118_AQ),
.I3(CLBLM_L_X94Y124_SLICE_X148Y124_DO6),
.I4(CLBLM_L_X90Y117_SLICE_X143Y117_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y119_SLICE_X143Y119_DO5),
.O6(CLBLM_L_X90Y119_SLICE_X143Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_CLUT (
.I0(CLBLM_L_X90Y120_SLICE_X143Y120_CQ),
.I1(CLBLM_L_X90Y119_SLICE_X143Y119_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y119_SLICE_X142Y119_C5Q),
.I4(CLBLM_L_X90Y119_SLICE_X143Y119_B5Q),
.I5(CLBLM_L_X90Y120_SLICE_X143Y120_BQ),
.O5(CLBLM_L_X90Y119_SLICE_X143Y119_CO5),
.O6(CLBLM_L_X90Y119_SLICE_X143Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f000f000)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y120_SLICE_X143Y120_CQ),
.I4(CLBLM_R_X93Y124_SLICE_X147Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y119_SLICE_X143Y119_BO5),
.O6(CLBLM_L_X90Y119_SLICE_X143Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_L_X90Y119_SLICE_X143Y119_ALUT (
.I0(CLBLM_L_X90Y119_SLICE_X143Y119_B5Q),
.I1(CLBLM_L_X90Y120_SLICE_X143Y120_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y119_SLICE_X143Y119_CQ),
.I4(CLBLM_L_X90Y120_SLICE_X143Y120_CQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y119_SLICE_X143Y119_AO5),
.O6(CLBLM_L_X90Y119_SLICE_X143Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X142Y120_AO5),
.Q(CLBLM_L_X90Y120_SLICE_X142Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X142Y120_CO5),
.Q(CLBLM_L_X90Y120_SLICE_X142Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X142Y120_AO6),
.Q(CLBLM_L_X90Y120_SLICE_X142Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X142Y120_BO6),
.Q(CLBLM_L_X90Y120_SLICE_X142Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0069699696)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_DLUT (
.I0(CLBLM_L_X90Y120_SLICE_X142Y120_BQ),
.I1(CLBLM_R_X89Y120_SLICE_X141Y120_AQ),
.I2(CLBLM_L_X90Y120_SLICE_X143Y120_C5Q),
.I3(CLBLM_L_X90Y119_SLICE_X142Y119_CQ),
.I4(CLBLM_L_X90Y120_SLICE_X142Y120_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y120_SLICE_X142Y120_DO5),
.O6(CLBLM_L_X90Y120_SLICE_X142Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696f000f000)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_CLUT (
.I0(CLBLM_L_X90Y120_SLICE_X142Y120_BQ),
.I1(CLBLM_R_X89Y120_SLICE_X141Y120_AQ),
.I2(CLBLM_L_X90Y120_SLICE_X143Y120_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y120_SLICE_X142Y120_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y120_SLICE_X142Y120_CO5),
.O6(CLBLM_L_X90Y120_SLICE_X142Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e020e0e0202020)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_BLUT (
.I0(CLBLM_R_X93Y124_SLICE_X146Y124_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X90Y120_SLICE_X142Y120_A5Q),
.I5(CLBLM_L_X90Y120_SLICE_X142Y120_CO6),
.O5(CLBLM_L_X90Y120_SLICE_X142Y120_BO5),
.O6(CLBLM_L_X90Y120_SLICE_X142Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X90Y120_SLICE_X142Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y120_SLICE_X142Y120_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X89Y122_SLICE_X141Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y120_SLICE_X142Y120_AO5),
.O6(CLBLM_L_X90Y120_SLICE_X142Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X143Y120_AO5),
.Q(CLBLM_L_X90Y120_SLICE_X143Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X143Y120_CO5),
.Q(CLBLM_L_X90Y120_SLICE_X143Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X143Y120_AO6),
.Q(CLBLM_L_X90Y120_SLICE_X143Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X143Y120_BO6),
.Q(CLBLM_L_X90Y120_SLICE_X143Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y120_SLICE_X143Y120_CO6),
.Q(CLBLM_L_X90Y120_SLICE_X143Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y120_SLICE_X143Y120_DO5),
.O6(CLBLM_L_X90Y120_SLICE_X143Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y120_SLICE_X141Y120_AQ),
.I2(CLBLM_L_X90Y120_SLICE_X143Y120_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y120_SLICE_X143Y120_CO5),
.O6(CLBLM_L_X90Y120_SLICE_X143Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b07030c0804000)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y119_SLICE_X143Y119_AO6),
.I4(CLBLM_L_X90Y120_SLICE_X142Y120_AQ),
.I5(CLBLM_L_X94Y123_SLICE_X148Y123_DO6),
.O5(CLBLM_L_X90Y120_SLICE_X143Y120_BO5),
.O6(CLBLM_L_X90Y120_SLICE_X143Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222220aa0a00a)
  ) CLBLM_L_X90Y120_SLICE_X143Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y117_SLICE_X143Y117_CO6),
.I2(CLBLM_L_X92Y122_SLICE_X144Y122_C5Q),
.I3(CLBLM_L_X90Y116_SLICE_X143Y116_B5Q),
.I4(CLBLM_L_X90Y122_SLICE_X143Y122_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y120_SLICE_X143Y120_AO5),
.O6(CLBLM_L_X90Y120_SLICE_X143Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y121_SLICE_X142Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y121_SLICE_X142Y121_AO5),
.Q(CLBLM_L_X90Y121_SLICE_X142Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y121_SLICE_X142Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y121_SLICE_X142Y121_AO6),
.Q(CLBLM_L_X90Y121_SLICE_X142Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y121_SLICE_X142Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y121_SLICE_X142Y121_DO5),
.O6(CLBLM_L_X90Y121_SLICE_X142Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y121_SLICE_X142Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y121_SLICE_X142Y121_CO5),
.O6(CLBLM_L_X90Y121_SLICE_X142Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y121_SLICE_X142Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y121_SLICE_X142Y121_BO5),
.O6(CLBLM_L_X90Y121_SLICE_X142Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0a0a0a0a0)
  ) CLBLM_L_X90Y121_SLICE_X142Y121_ALUT (
.I0(CLBLM_L_X90Y114_SLICE_X142Y114_A5Q),
.I1(CLBLM_L_X90Y121_SLICE_X142Y121_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y121_SLICE_X142Y121_AO5),
.O6(CLBLM_L_X90Y121_SLICE_X142Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y121_SLICE_X143Y121_BO5),
.Q(CLBLM_L_X90Y121_SLICE_X143Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y121_SLICE_X143Y121_CO5),
.Q(CLBLM_L_X90Y121_SLICE_X143Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y121_SLICE_X143Y121_AO6),
.Q(CLBLM_L_X90Y121_SLICE_X143Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y121_SLICE_X143Y121_CO6),
.Q(CLBLM_L_X90Y121_SLICE_X143Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_DLUT (
.I0(CLBLM_L_X90Y121_SLICE_X143Y121_C5Q),
.I1(CLBLM_L_X90Y121_SLICE_X143Y121_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y121_SLICE_X143Y121_A5Q),
.I4(CLBLM_L_X90Y121_SLICE_X143Y121_AQ),
.I5(CLBLM_L_X92Y121_SLICE_X145Y121_CQ),
.O5(CLBLM_L_X90Y121_SLICE_X143Y121_DO5),
.O6(CLBLM_L_X90Y121_SLICE_X143Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y121_SLICE_X143Y121_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X90Y121_SLICE_X143Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y121_SLICE_X143Y121_CO5),
.O6(CLBLM_L_X90Y121_SLICE_X143Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_BLUT (
.I0(CLBLM_L_X90Y121_SLICE_X143Y121_AQ),
.I1(CLBLM_L_X90Y121_SLICE_X143Y121_A5Q),
.I2(CLBLM_L_X90Y121_SLICE_X143Y121_CQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y121_SLICE_X143Y121_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y121_SLICE_X143Y121_BO5),
.O6(CLBLM_L_X90Y121_SLICE_X143Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e20000ee220000)
  ) CLBLM_L_X90Y121_SLICE_X143Y121_ALUT (
.I0(CLBLM_R_X89Y125_SLICE_X141Y125_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X90Y121_SLICE_X142Y121_A5Q),
.I3(CLBLM_L_X90Y121_SLICE_X143Y121_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y121_SLICE_X143Y121_AO5),
.O6(CLBLM_L_X90Y121_SLICE_X143Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X142Y122_AO5),
.Q(CLBLM_L_X90Y122_SLICE_X142Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X142Y122_AO6),
.Q(CLBLM_L_X90Y122_SLICE_X142Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X142Y122_BO6),
.Q(CLBLM_L_X90Y122_SLICE_X142Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y122_SLICE_X142Y122_DO5),
.O6(CLBLM_L_X90Y122_SLICE_X142Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y122_SLICE_X142Y122_CO5),
.O6(CLBLM_L_X90Y122_SLICE_X142Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c000c0a0a0a0a0)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_BLUT (
.I0(CLBLM_L_X90Y128_SLICE_X142Y128_DO6),
.I1(CLBLM_L_X92Y122_SLICE_X144Y122_AO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X90Y122_SLICE_X142Y122_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X90Y122_SLICE_X142Y122_BO5),
.O6(CLBLM_L_X90Y122_SLICE_X142Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_L_X90Y122_SLICE_X142Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y122_SLICE_X142Y122_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y121_SLICE_X142Y121_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y122_SLICE_X142Y122_AO5),
.O6(CLBLM_L_X90Y122_SLICE_X142Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X143Y122_BO5),
.Q(CLBLM_L_X90Y122_SLICE_X143Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X143Y122_CO5),
.Q(CLBLM_L_X90Y122_SLICE_X143Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X143Y122_AO6),
.Q(CLBLM_L_X90Y122_SLICE_X143Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y122_SLICE_X143Y122_CO6),
.Q(CLBLM_L_X90Y122_SLICE_X143Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_DLUT (
.I0(CLBLM_R_X89Y120_SLICE_X141Y120_BQ),
.I1(CLBLM_L_X90Y122_SLICE_X143Y122_CQ),
.I2(CLBLM_L_X90Y124_SLICE_X143Y124_B5Q),
.I3(CLBLM_L_X90Y122_SLICE_X143Y122_A5Q),
.I4(CLBLM_L_X90Y122_SLICE_X143Y122_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y122_SLICE_X143Y122_DO5),
.O6(CLBLM_L_X90Y122_SLICE_X143Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aa00aa00)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X92Y120_SLICE_X144Y120_B5Q),
.I4(CLBLM_L_X90Y122_SLICE_X143Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y122_SLICE_X143Y122_CO5),
.O6(CLBLM_L_X90Y122_SLICE_X143Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966c0c0c0c0)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_BLUT (
.I0(CLBLM_L_X90Y122_SLICE_X143Y122_AQ),
.I1(CLBLM_L_X90Y124_SLICE_X143Y124_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y122_SLICE_X143Y122_CQ),
.I4(CLBLM_L_X90Y122_SLICE_X143Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y122_SLICE_X143Y122_BO5),
.O6(CLBLM_L_X90Y122_SLICE_X143Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0e0202020e020)
  ) CLBLM_L_X90Y122_SLICE_X143Y122_ALUT (
.I0(CLBLM_R_X93Y128_SLICE_X146Y128_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y122_SLICE_X143Y122_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y124_SLICE_X141Y124_AQ),
.O5(CLBLM_L_X90Y122_SLICE_X143Y122_AO5),
.O6(CLBLM_L_X90Y122_SLICE_X143Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X142Y123_AO5),
.Q(CLBLM_L_X90Y123_SLICE_X142Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X142Y123_BO5),
.Q(CLBLM_L_X90Y123_SLICE_X142Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X142Y123_CO5),
.Q(CLBLM_L_X90Y123_SLICE_X142Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X142Y123_AO6),
.Q(CLBLM_L_X90Y123_SLICE_X142Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X142Y123_BO6),
.Q(CLBLM_L_X90Y123_SLICE_X142Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X142Y123_CO6),
.Q(CLBLM_L_X90Y123_SLICE_X142Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y123_SLICE_X142Y123_DO5),
.O6(CLBLM_L_X90Y123_SLICE_X142Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00aa00a88882222)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y124_SLICE_X142Y124_A5Q),
.I2(CLBLM_R_X89Y123_SLICE_X141Y123_A5Q),
.I3(CLBLM_L_X92Y122_SLICE_X144Y122_AQ),
.I4(CLBLM_L_X90Y123_SLICE_X142Y123_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y123_SLICE_X142Y123_CO5),
.O6(CLBLM_L_X90Y123_SLICE_X142Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0303060906090)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_BLUT (
.I0(CLBLM_L_X90Y123_SLICE_X142Y123_CQ),
.I1(CLBLM_L_X90Y115_SLICE_X142Y115_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y123_SLICE_X143Y123_A5Q),
.I4(CLBLM_L_X92Y121_SLICE_X145Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y123_SLICE_X142Y123_BO5),
.O6(CLBLM_L_X90Y123_SLICE_X142Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0a0a0a0a0)
  ) CLBLM_L_X90Y123_SLICE_X142Y123_ALUT (
.I0(CLBLM_L_X90Y122_SLICE_X142Y122_AQ),
.I1(CLBLM_L_X90Y123_SLICE_X142Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y123_SLICE_X142Y123_AO5),
.O6(CLBLM_L_X90Y123_SLICE_X142Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X143Y123_BO5),
.Q(CLBLM_L_X90Y123_SLICE_X143Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X143Y123_CO5),
.Q(CLBLM_L_X90Y123_SLICE_X143Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X143Y123_AO6),
.Q(CLBLM_L_X90Y123_SLICE_X143Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y123_SLICE_X143Y123_CO6),
.Q(CLBLM_L_X90Y123_SLICE_X143Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_DLUT (
.I0(CLBLM_L_X90Y123_SLICE_X143Y123_C5Q),
.I1(CLBLM_L_X90Y123_SLICE_X143Y123_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y123_SLICE_X143Y123_A5Q),
.I4(CLBLM_L_X90Y123_SLICE_X143Y123_AQ),
.I5(CLBLM_L_X92Y121_SLICE_X144Y121_D5Q),
.O5(CLBLM_L_X90Y123_SLICE_X143Y123_DO5),
.O6(CLBLM_L_X90Y123_SLICE_X143Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y123_SLICE_X143Y123_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X90Y123_SLICE_X143Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y123_SLICE_X143Y123_CO5),
.O6(CLBLM_L_X90Y123_SLICE_X143Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_BLUT (
.I0(CLBLM_L_X90Y123_SLICE_X143Y123_AQ),
.I1(CLBLM_L_X90Y123_SLICE_X143Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y123_SLICE_X143Y123_CQ),
.I4(CLBLM_L_X90Y123_SLICE_X143Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y123_SLICE_X143Y123_BO5),
.O6(CLBLM_L_X90Y123_SLICE_X143Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b0f0308080c000)
  ) CLBLM_L_X90Y123_SLICE_X143Y123_ALUT (
.I0(CLBLM_L_X90Y122_SLICE_X142Y122_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y123_SLICE_X143Y123_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X90Y124_SLICE_X143Y124_DO6),
.O5(CLBLM_L_X90Y123_SLICE_X143Y123_AO5),
.O6(CLBLM_L_X90Y123_SLICE_X143Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X142Y124_BO5),
.Q(CLBLM_L_X90Y124_SLICE_X142Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X142Y124_CO5),
.Q(CLBLM_L_X90Y124_SLICE_X142Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X142Y124_AO6),
.Q(CLBLM_L_X90Y124_SLICE_X142Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X142Y124_CO6),
.Q(CLBLM_L_X90Y124_SLICE_X142Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_DLUT (
.I0(CLBLM_L_X90Y124_SLICE_X142Y124_C5Q),
.I1(CLBLM_L_X90Y124_SLICE_X142Y124_CQ),
.I2(CLBLM_L_X90Y124_SLICE_X142Y124_AQ),
.I3(CLBLM_L_X90Y124_SLICE_X142Y124_A5Q),
.I4(CLBLM_L_X92Y122_SLICE_X145Y122_C5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y124_SLICE_X142Y124_DO5),
.O6(CLBLM_L_X90Y124_SLICE_X142Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y124_SLICE_X142Y124_CQ),
.I2(CLBLM_L_X90Y124_SLICE_X142Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y124_SLICE_X142Y124_CO5),
.O6(CLBLM_L_X90Y124_SLICE_X142Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_BLUT (
.I0(CLBLM_L_X90Y124_SLICE_X142Y124_AQ),
.I1(CLBLM_L_X90Y124_SLICE_X142Y124_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y124_SLICE_X142Y124_CQ),
.I4(CLBLM_L_X90Y124_SLICE_X142Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y124_SLICE_X142Y124_BO5),
.O6(CLBLM_L_X90Y124_SLICE_X142Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e02020e020e020)
  ) CLBLM_L_X90Y124_SLICE_X142Y124_ALUT (
.I0(CLBLM_L_X90Y128_SLICE_X142Y128_CO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y124_SLICE_X142Y124_BO6),
.I4(CLBLM_L_X90Y123_SLICE_X142Y123_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y124_SLICE_X142Y124_AO5),
.O6(CLBLM_L_X90Y124_SLICE_X142Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X143Y124_BO5),
.Q(CLBLM_L_X90Y124_SLICE_X143Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X143Y124_CO5),
.Q(CLBLM_L_X90Y124_SLICE_X143Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X143Y124_AO5),
.Q(CLBLM_L_X90Y124_SLICE_X143Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X143Y124_BO6),
.Q(CLBLM_L_X90Y124_SLICE_X143Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y124_SLICE_X143Y124_CO6),
.Q(CLBLM_L_X90Y124_SLICE_X143Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_DLUT (
.I0(CLBLM_L_X90Y124_SLICE_X143Y124_BQ),
.I1(CLBLM_L_X90Y124_SLICE_X143Y124_AQ),
.I2(CLBLM_L_X90Y123_SLICE_X142Y123_B5Q),
.I3(CLBLM_L_X90Y125_SLICE_X142Y125_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X90Y128_SLICE_X143Y128_BQ),
.O5(CLBLM_L_X90Y124_SLICE_X143Y124_DO5),
.O6(CLBLM_L_X90Y124_SLICE_X143Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0000aa82828282)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y124_SLICE_X143Y124_CQ),
.I2(CLBLM_R_X89Y121_SLICE_X141Y121_A5Q),
.I3(CLBLM_R_X89Y122_SLICE_X141Y122_B5Q),
.I4(CLBLM_L_X90Y125_SLICE_X143Y125_DQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y124_SLICE_X143Y124_CO5),
.O6(CLBLM_L_X90Y124_SLICE_X143Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y122_SLICE_X143Y122_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y128_SLICE_X143Y128_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y124_SLICE_X143Y124_BO5),
.O6(CLBLM_L_X90Y124_SLICE_X143Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_L_X90Y124_SLICE_X143Y124_ALUT (
.I0(CLBLM_L_X90Y125_SLICE_X142Y125_A5Q),
.I1(CLBLM_L_X90Y128_SLICE_X143Y128_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y124_SLICE_X143Y124_AQ),
.I4(CLBLM_L_X90Y124_SLICE_X143Y124_BQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y124_SLICE_X143Y124_AO5),
.O6(CLBLM_L_X90Y124_SLICE_X143Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X142Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X142Y125_AO5),
.Q(CLBLM_L_X90Y125_SLICE_X142Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X142Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X142Y125_AO6),
.Q(CLBLM_L_X90Y125_SLICE_X142Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y125_SLICE_X142Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y125_SLICE_X142Y125_DO5),
.O6(CLBLM_L_X90Y125_SLICE_X142Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y125_SLICE_X142Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y125_SLICE_X142Y125_CO5),
.O6(CLBLM_L_X90Y125_SLICE_X142Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd8d88dd88d8dd8)
  ) CLBLM_L_X90Y125_SLICE_X142Y125_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X90Y123_SLICE_X142Y123_BQ),
.I2(CLBLM_L_X90Y125_SLICE_X142Y125_AQ),
.I3(CLBLM_R_X89Y125_SLICE_X141Y125_C5Q),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_BQ),
.I5(CLBLM_R_X89Y125_SLICE_X140Y125_B5Q),
.O5(CLBLM_L_X90Y125_SLICE_X142Y125_BO5),
.O6(CLBLM_L_X90Y125_SLICE_X142Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f000f000)
  ) CLBLM_L_X90Y125_SLICE_X142Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y124_SLICE_X143Y124_BQ),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_BQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y125_SLICE_X142Y125_AO5),
.O6(CLBLM_L_X90Y125_SLICE_X142Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X143Y125_AO5),
.Q(CLBLM_L_X90Y125_SLICE_X143Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X143Y125_BO5),
.Q(CLBLM_L_X90Y125_SLICE_X143Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X143Y125_AO6),
.Q(CLBLM_L_X90Y125_SLICE_X143Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X143Y125_BO6),
.Q(CLBLM_L_X90Y125_SLICE_X143Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X143Y125_CO6),
.Q(CLBLM_L_X90Y125_SLICE_X143Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y125_SLICE_X143Y125_DO6),
.Q(CLBLM_L_X90Y125_SLICE_X143Y125_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222888888882222)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y125_SLICE_X143Y125_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X90Y116_SLICE_X143Y116_B5Q),
.I5(CLBLM_L_X90Y122_SLICE_X143Y122_A5Q),
.O5(CLBLM_L_X90Y125_SLICE_X143Y125_DO5),
.O6(CLBLM_L_X90Y125_SLICE_X143Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a00a0a0a0a)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X92Y131_SLICE_X144Y131_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X89Y124_SLICE_X140Y124_BQ),
.O5(CLBLM_L_X90Y125_SLICE_X143Y125_CO5),
.O6(CLBLM_L_X90Y125_SLICE_X143Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha050a05060609090)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_BLUT (
.I0(CLBLM_L_X90Y116_SLICE_X143Y116_B5Q),
.I1(CLBLM_L_X90Y124_SLICE_X143Y124_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y125_SLICE_X140Y125_B5Q),
.I4(CLBLM_L_X90Y128_SLICE_X143Y128_DQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y125_SLICE_X143Y125_BO5),
.O6(CLBLM_L_X90Y125_SLICE_X143Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X90Y125_SLICE_X143Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y125_SLICE_X143Y125_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y123_SLICE_X142Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y125_SLICE_X143Y125_AO5),
.O6(CLBLM_L_X90Y125_SLICE_X143Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X142Y126_BO5),
.Q(CLBLM_L_X90Y126_SLICE_X142Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X142Y126_CO5),
.Q(CLBLM_L_X90Y126_SLICE_X142Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X142Y126_AO5),
.Q(CLBLM_L_X90Y126_SLICE_X142Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X142Y126_BO6),
.Q(CLBLM_L_X90Y126_SLICE_X142Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X142Y126_CO6),
.Q(CLBLM_L_X90Y126_SLICE_X142Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_DLUT (
.I0(CLBLM_L_X90Y126_SLICE_X142Y126_BQ),
.I1(CLBLM_L_X90Y126_SLICE_X142Y126_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y123_SLICE_X144Y123_DQ),
.I4(CLBLM_L_X90Y126_SLICE_X142Y126_B5Q),
.I5(CLBLM_R_X89Y126_SLICE_X140Y126_AQ),
.O5(CLBLM_L_X90Y126_SLICE_X142Y126_DO5),
.O6(CLBLM_L_X90Y126_SLICE_X142Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_CLUT (
.I0(CLBLM_L_X90Y126_SLICE_X142Y126_CQ),
.I1(CLBLM_L_X90Y126_SLICE_X143Y126_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y124_SLICE_X144Y124_A5Q),
.I4(CLBLM_L_X90Y123_SLICE_X142Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y126_SLICE_X142Y126_CO5),
.O6(CLBLM_L_X90Y126_SLICE_X142Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y126_SLICE_X142Y126_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y126_SLICE_X140Y126_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y126_SLICE_X142Y126_BO5),
.O6(CLBLM_L_X90Y126_SLICE_X142Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_L_X90Y126_SLICE_X142Y126_ALUT (
.I0(CLBLM_L_X90Y126_SLICE_X142Y126_B5Q),
.I1(CLBLM_L_X90Y126_SLICE_X142Y126_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y126_SLICE_X140Y126_AQ),
.I4(CLBLM_L_X90Y126_SLICE_X142Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y126_SLICE_X142Y126_AO5),
.O6(CLBLM_L_X90Y126_SLICE_X142Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X143Y126_BO5),
.Q(CLBLM_L_X90Y126_SLICE_X143Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X143Y126_CO5),
.Q(CLBLM_L_X90Y126_SLICE_X143Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X143Y126_AO6),
.Q(CLBLM_L_X90Y126_SLICE_X143Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y126_SLICE_X143Y126_CO6),
.Q(CLBLM_L_X90Y126_SLICE_X143Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cacac5cac5c5ca)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_DLUT (
.I0(CLBLM_L_X90Y126_SLICE_X143Y126_C5Q),
.I1(CLBLM_L_X92Y124_SLICE_X145Y124_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y126_SLICE_X143Y126_A5Q),
.I4(CLBLM_L_X90Y126_SLICE_X143Y126_AQ),
.I5(CLBLM_L_X90Y126_SLICE_X143Y126_CQ),
.O5(CLBLM_L_X90Y126_SLICE_X143Y126_DO5),
.O6(CLBLM_L_X90Y126_SLICE_X143Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y126_SLICE_X143Y126_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X90Y126_SLICE_X143Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y126_SLICE_X143Y126_CO5),
.O6(CLBLM_L_X90Y126_SLICE_X143Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_BLUT (
.I0(CLBLM_L_X90Y126_SLICE_X143Y126_AQ),
.I1(CLBLM_L_X90Y126_SLICE_X143Y126_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y126_SLICE_X143Y126_CQ),
.I4(CLBLM_L_X90Y126_SLICE_X143Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y126_SLICE_X143Y126_BO5),
.O6(CLBLM_L_X90Y126_SLICE_X143Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c03000a0a0a0a0)
  ) CLBLM_L_X90Y126_SLICE_X143Y126_ALUT (
.I0(CLBLM_L_X90Y131_SLICE_X142Y131_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y126_SLICE_X143Y126_BO6),
.I4(CLBLM_L_X90Y125_SLICE_X143Y125_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X90Y126_SLICE_X143Y126_AO5),
.O6(CLBLM_L_X90Y126_SLICE_X143Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X142Y128_BO5),
.Q(CLBLM_L_X90Y128_SLICE_X142Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X142Y128_AO5),
.Q(CLBLM_L_X90Y128_SLICE_X142Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X142Y128_BO6),
.Q(CLBLM_L_X90Y128_SLICE_X142Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_DLUT (
.I0(CLBLM_L_X90Y123_SLICE_X142Y123_CQ),
.I1(CLBLM_L_X90Y128_SLICE_X142Y128_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y128_SLICE_X143Y128_CQ),
.I4(CLBLM_L_X90Y128_SLICE_X142Y128_B5Q),
.I5(CLBLM_R_X89Y128_SLICE_X141Y128_AQ),
.O5(CLBLM_L_X90Y128_SLICE_X142Y128_DO5),
.O6(CLBLM_L_X90Y128_SLICE_X142Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_CLUT (
.I0(CLBLM_L_X90Y129_SLICE_X142Y129_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X90Y128_SLICE_X142Y128_BQ),
.I3(CLBLM_L_X90Y129_SLICE_X142Y129_C5Q),
.I4(CLBLM_L_X90Y129_SLICE_X142Y129_A5Q),
.I5(CLBLM_L_X90Y123_SLICE_X142Y123_C5Q),
.O5(CLBLM_L_X90Y128_SLICE_X142Y128_CO5),
.O6(CLBLM_L_X90Y128_SLICE_X142Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f000f000)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y128_SLICE_X141Y128_AQ),
.I4(CLBLM_L_X90Y129_SLICE_X142Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y128_SLICE_X142Y128_BO5),
.O6(CLBLM_L_X90Y128_SLICE_X142Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_L_X90Y128_SLICE_X142Y128_ALUT (
.I0(CLBLM_L_X90Y128_SLICE_X142Y128_B5Q),
.I1(CLBLM_L_X90Y128_SLICE_X142Y128_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y128_SLICE_X141Y128_AQ),
.I4(CLBLM_L_X90Y128_SLICE_X143Y128_CQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y128_SLICE_X142Y128_AO5),
.O6(CLBLM_L_X90Y128_SLICE_X142Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X143Y128_AO5),
.Q(CLBLM_L_X90Y128_SLICE_X143Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X143Y128_DO5),
.Q(CLBLM_L_X90Y128_SLICE_X143Y128_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X143Y128_AO6),
.Q(CLBLM_L_X90Y128_SLICE_X143Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X143Y128_BO6),
.Q(CLBLM_L_X90Y128_SLICE_X143Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X143Y128_CO6),
.Q(CLBLM_L_X90Y128_SLICE_X143Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y128_SLICE_X143Y128_DO6),
.Q(CLBLM_L_X90Y128_SLICE_X143Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa550000c3c30000)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_DLUT (
.I0(CLBLM_L_X90Y128_SLICE_X142Y128_AQ),
.I1(CLBLM_L_X90Y125_SLICE_X143Y125_B5Q),
.I2(CLBLM_L_X90Y129_SLICE_X142Y129_A5Q),
.I3(CLBLM_L_X92Y126_SLICE_X145Y126_C5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y128_SLICE_X143Y128_DO5),
.O6(CLBLM_L_X90Y128_SLICE_X143Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e40000ff000000)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X90Y128_SLICE_X142Y128_AO6),
.I2(CLBLM_R_X89Y127_SLICE_X141Y127_AQ),
.I3(CLBLM_L_X92Y129_SLICE_X145Y129_DO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X90Y128_SLICE_X143Y128_CO5),
.O6(CLBLM_L_X90Y128_SLICE_X143Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0c0c000a0c0c0)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_BLUT (
.I0(CLBLM_L_X90Y124_SLICE_X143Y124_AO6),
.I1(CLBLM_L_X92Y128_SLICE_X145Y128_DO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X90Y128_SLICE_X143Y128_A5Q),
.O5(CLBLM_L_X90Y128_SLICE_X143Y128_BO5),
.O6(CLBLM_L_X90Y128_SLICE_X143Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X90Y128_SLICE_X143Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X90Y128_SLICE_X143Y128_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X89Y127_SLICE_X141Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X90Y128_SLICE_X143Y128_AO5),
.O6(CLBLM_L_X90Y128_SLICE_X143Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y129_SLICE_X142Y129_BO5),
.Q(CLBLM_L_X90Y129_SLICE_X142Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y129_SLICE_X142Y129_CO5),
.Q(CLBLM_L_X90Y129_SLICE_X142Y129_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y129_SLICE_X142Y129_AO6),
.Q(CLBLM_L_X90Y129_SLICE_X142Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y129_SLICE_X142Y129_CO6),
.Q(CLBLM_L_X90Y129_SLICE_X142Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X142Y129_DO5),
.O6(CLBLM_L_X90Y129_SLICE_X142Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X90Y130_SLICE_X142Y130_BQ),
.I3(CLBLM_L_X90Y128_SLICE_X142Y128_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X142Y129_CO5),
.O6(CLBLM_L_X90Y129_SLICE_X142Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_BLUT (
.I0(CLBLM_L_X90Y129_SLICE_X142Y129_AQ),
.I1(CLBLM_L_X90Y129_SLICE_X142Y129_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y128_SLICE_X142Y128_BQ),
.I4(CLBLM_L_X90Y129_SLICE_X142Y129_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X142Y129_BO5),
.O6(CLBLM_L_X90Y129_SLICE_X142Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0a0a0f000a0a0)
  ) CLBLM_L_X90Y129_SLICE_X142Y129_ALUT (
.I0(CLBLM_R_X93Y131_SLICE_X146Y131_DO6),
.I1(CLBLM_L_X90Y128_SLICE_X143Y128_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y129_SLICE_X142Y129_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y129_SLICE_X142Y129_AO5),
.O6(CLBLM_L_X90Y129_SLICE_X142Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y129_SLICE_X143Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X143Y129_DO5),
.O6(CLBLM_L_X90Y129_SLICE_X143Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y129_SLICE_X143Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X143Y129_CO5),
.O6(CLBLM_L_X90Y129_SLICE_X143Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y129_SLICE_X143Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X143Y129_BO5),
.O6(CLBLM_L_X90Y129_SLICE_X143Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y129_SLICE_X143Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y129_SLICE_X143Y129_AO5),
.O6(CLBLM_L_X90Y129_SLICE_X143Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y130_SLICE_X142Y130_AO5),
.Q(CLBLM_L_X90Y130_SLICE_X142Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y130_SLICE_X142Y130_CO5),
.Q(CLBLM_L_X90Y130_SLICE_X142Y130_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y130_SLICE_X142Y130_AO6),
.Q(CLBLM_L_X90Y130_SLICE_X142Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y130_SLICE_X142Y130_BO6),
.Q(CLBLM_L_X90Y130_SLICE_X142Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_DLUT (
.I0(CLBLM_L_X90Y131_SLICE_X142Y131_C5Q),
.I1(CLBLM_L_X90Y126_SLICE_X142Y126_CQ),
.I2(CLBLM_L_X90Y129_SLICE_X142Y129_CQ),
.I3(CLBLM_L_X90Y130_SLICE_X142Y130_BQ),
.I4(CLBLM_L_X90Y130_SLICE_X142Y130_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y130_SLICE_X142Y130_DO5),
.O6(CLBLM_L_X90Y130_SLICE_X142Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996aaaa0000)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_CLUT (
.I0(CLBLM_L_X90Y131_SLICE_X142Y131_C5Q),
.I1(CLBLM_L_X90Y130_SLICE_X142Y130_B5Q),
.I2(CLBLM_L_X90Y129_SLICE_X142Y129_CQ),
.I3(CLBLM_L_X90Y130_SLICE_X142Y130_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y130_SLICE_X142Y130_CO5),
.O6(CLBLM_L_X90Y130_SLICE_X142Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88aaa0a08800a0a0)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y130_SLICE_X142Y130_A5Q),
.I2(CLBLM_L_X92Y131_SLICE_X144Y131_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X90Y130_SLICE_X142Y130_CO6),
.O5(CLBLM_L_X90Y130_SLICE_X142Y130_BO5),
.O6(CLBLM_L_X90Y130_SLICE_X142Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X90Y130_SLICE_X142Y130_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y130_SLICE_X142Y130_A5Q),
.I2(CLBLM_L_X90Y128_SLICE_X143Y128_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y130_SLICE_X142Y130_AO5),
.O6(CLBLM_L_X90Y130_SLICE_X142Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y130_SLICE_X143Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y130_SLICE_X143Y130_DO5),
.O6(CLBLM_L_X90Y130_SLICE_X143Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y130_SLICE_X143Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y130_SLICE_X143Y130_CO5),
.O6(CLBLM_L_X90Y130_SLICE_X143Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y130_SLICE_X143Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y130_SLICE_X143Y130_BO5),
.O6(CLBLM_L_X90Y130_SLICE_X143Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y130_SLICE_X143Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y130_SLICE_X143Y130_AO5),
.O6(CLBLM_L_X90Y130_SLICE_X143Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y131_SLICE_X142Y131_BO5),
.Q(CLBLM_L_X90Y131_SLICE_X142Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y131_SLICE_X142Y131_CO5),
.Q(CLBLM_L_X90Y131_SLICE_X142Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y131_SLICE_X142Y131_AO6),
.Q(CLBLM_L_X90Y131_SLICE_X142Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X90Y131_SLICE_X142Y131_CO6),
.Q(CLBLM_L_X90Y131_SLICE_X142Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_DLUT (
.I0(CLBLM_L_X90Y126_SLICE_X142Y126_C5Q),
.I1(CLBLM_L_X90Y131_SLICE_X142Y131_CQ),
.I2(CLBLM_L_X90Y131_SLICE_X142Y131_AQ),
.I3(CLBLM_L_X90Y131_SLICE_X142Y131_A5Q),
.I4(CLBLM_R_X89Y131_SLICE_X140Y131_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X90Y131_SLICE_X142Y131_DO5),
.O6(CLBLM_L_X90Y131_SLICE_X142Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y131_SLICE_X142Y131_AQ),
.I2(1'b1),
.I3(CLBLM_L_X90Y129_SLICE_X142Y129_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y131_SLICE_X142Y131_CO5),
.O6(CLBLM_L_X90Y131_SLICE_X142Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996aaaa0000)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_BLUT (
.I0(CLBLM_R_X89Y131_SLICE_X140Y131_A5Q),
.I1(CLBLM_L_X90Y131_SLICE_X142Y131_A5Q),
.I2(CLBLM_L_X90Y131_SLICE_X142Y131_AQ),
.I3(CLBLM_L_X90Y131_SLICE_X142Y131_CQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X90Y131_SLICE_X142Y131_BO5),
.O6(CLBLM_L_X90Y131_SLICE_X142Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc00000aaaa0000)
  ) CLBLM_L_X90Y131_SLICE_X142Y131_ALUT (
.I0(CLBLM_R_X93Y133_SLICE_X146Y133_DO6),
.I1(CLBLM_L_X90Y130_SLICE_X142Y130_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X90Y131_SLICE_X142Y131_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X90Y131_SLICE_X142Y131_AO5),
.O6(CLBLM_L_X90Y131_SLICE_X142Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y131_SLICE_X143Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y131_SLICE_X143Y131_DO5),
.O6(CLBLM_L_X90Y131_SLICE_X143Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y131_SLICE_X143Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y131_SLICE_X143Y131_CO5),
.O6(CLBLM_L_X90Y131_SLICE_X143Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y131_SLICE_X143Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y131_SLICE_X143Y131_BO5),
.O6(CLBLM_L_X90Y131_SLICE_X143Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X90Y131_SLICE_X143Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X90Y131_SLICE_X143Y131_AO5),
.O6(CLBLM_L_X90Y131_SLICE_X143Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y112_SLICE_X144Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X144Y112_DO5),
.O6(CLBLM_L_X92Y112_SLICE_X144Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y112_SLICE_X144Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X144Y112_CO5),
.O6(CLBLM_L_X92Y112_SLICE_X144Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y112_SLICE_X144Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X144Y112_BO5),
.O6(CLBLM_L_X92Y112_SLICE_X144Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y112_SLICE_X144Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X144Y112_AO5),
.O6(CLBLM_L_X92Y112_SLICE_X144Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y112_SLICE_X145Y112_AO5),
.Q(CLBLM_L_X92Y112_SLICE_X145Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y112_SLICE_X145Y112_BO5),
.Q(CLBLM_L_X92Y112_SLICE_X145Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y112_SLICE_X145Y112_AO6),
.Q(CLBLM_L_X92Y112_SLICE_X145Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y112_SLICE_X145Y112_BO6),
.Q(CLBLM_L_X92Y112_SLICE_X145Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X145Y112_DO5),
.O6(CLBLM_L_X92Y112_SLICE_X145Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X92Y112_SLICE_X145Y112_AQ),
.I2(1'b1),
.I3(CLBLM_L_X92Y112_SLICE_X145Y112_BQ),
.I4(CLBLM_L_X92Y112_SLICE_X145Y112_B5Q),
.I5(CLBLM_R_X93Y115_SLICE_X146Y115_AQ),
.O5(CLBLM_L_X92Y112_SLICE_X145Y112_CO5),
.O6(CLBLM_L_X92Y112_SLICE_X145Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y112_SLICE_X145Y112_AQ),
.I3(1'b1),
.I4(CLBLM_L_X92Y112_SLICE_X145Y112_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X145Y112_BO5),
.O6(CLBLM_L_X92Y112_SLICE_X145Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_L_X92Y112_SLICE_X145Y112_ALUT (
.I0(CLBLM_R_X93Y112_SLICE_X146Y112_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y115_SLICE_X146Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y112_SLICE_X145Y112_AO5),
.O6(CLBLM_L_X92Y112_SLICE_X145Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X144Y113_AO5),
.Q(CLBLM_L_X92Y113_SLICE_X144Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X144Y113_BO5),
.Q(CLBLM_L_X92Y113_SLICE_X144Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X144Y113_AO6),
.Q(CLBLM_L_X92Y113_SLICE_X144Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X144Y113_BO6),
.Q(CLBLM_L_X92Y113_SLICE_X144Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y113_SLICE_X144Y113_DO5),
.O6(CLBLM_L_X92Y113_SLICE_X144Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_CLUT (
.I0(CLBLM_L_X92Y113_SLICE_X145Y113_AQ),
.I1(CLBLM_L_X92Y113_SLICE_X144Y113_AQ),
.I2(CLBLM_L_X92Y113_SLICE_X144Y113_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X92Y113_SLICE_X144Y113_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y113_SLICE_X144Y113_CO5),
.O6(CLBLM_L_X92Y113_SLICE_X144Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y113_SLICE_X144Y113_AQ),
.I3(1'b1),
.I4(CLBLM_L_X92Y113_SLICE_X144Y113_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y113_SLICE_X144Y113_BO5),
.O6(CLBLM_L_X92Y113_SLICE_X144Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_L_X92Y113_SLICE_X144Y113_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y113_SLICE_X146Y113_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X92Y113_SLICE_X145Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y113_SLICE_X144Y113_AO5),
.O6(CLBLM_L_X92Y113_SLICE_X144Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X145Y113_AO5),
.Q(CLBLM_L_X92Y113_SLICE_X145Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X145Y113_BO5),
.Q(CLBLM_L_X92Y113_SLICE_X145Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X145Y113_AO6),
.Q(CLBLM_L_X92Y113_SLICE_X145Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y113_SLICE_X145Y113_BO6),
.Q(CLBLM_L_X92Y113_SLICE_X145Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5404f4a45e0efeae)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X93Y118_SLICE_X147Y118_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y112_SLICE_X146Y112_DO6),
.I4(CLBLM_L_X92Y113_SLICE_X145Y113_B5Q),
.I5(CLBLM_R_X93Y113_SLICE_X146Y113_A5Q),
.O5(CLBLM_L_X92Y113_SLICE_X145Y113_DO5),
.O6(CLBLM_L_X92Y113_SLICE_X145Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505ffcfc505f0c0c)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_CLUT (
.I0(CLBLM_L_X92Y113_SLICE_X145Y113_BQ),
.I1(CLBLM_L_X94Y116_SLICE_X148Y116_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X92Y113_SLICE_X145Y113_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X92Y112_SLICE_X145Y112_CO6),
.O5(CLBLM_L_X92Y113_SLICE_X145Y113_CO5),
.O6(CLBLM_L_X92Y113_SLICE_X145Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000cccc0000)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_BLUT (
.I0(CLBLM_L_X92Y113_SLICE_X145Y113_B5Q),
.I1(CLBLM_L_X94Y113_SLICE_X148Y113_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X92Y113_SLICE_X145Y113_BO5),
.O6(CLBLM_L_X92Y113_SLICE_X145Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500c300c300)
  ) CLBLM_L_X92Y113_SLICE_X145Y113_ALUT (
.I0(CLBLM_R_X93Y114_SLICE_X146Y114_CO6),
.I1(CLBLM_R_X93Y113_SLICE_X146Y113_A5Q),
.I2(CLBLM_L_X92Y112_SLICE_X145Y112_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y113_SLICE_X145Y113_AO5),
.O6(CLBLM_L_X92Y113_SLICE_X145Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y114_SLICE_X144Y114_AO5),
.Q(CLBLM_L_X92Y114_SLICE_X144Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y114_SLICE_X144Y114_BO5),
.Q(CLBLM_L_X92Y114_SLICE_X144Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y114_SLICE_X144Y114_AO6),
.Q(CLBLM_L_X92Y114_SLICE_X144Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y114_SLICE_X144Y114_BO6),
.Q(CLBLM_L_X92Y114_SLICE_X144Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_DLUT (
.I0(CLBLM_L_X90Y113_SLICE_X143Y113_BQ),
.I1(CLBLM_R_X93Y114_SLICE_X146Y114_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X92Y114_SLICE_X144Y114_BQ),
.I4(CLBLM_L_X92Y114_SLICE_X144Y114_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X144Y114_DO5),
.O6(CLBLM_L_X92Y114_SLICE_X144Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505f505ffcfc0c0c)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_CLUT (
.I0(CLBLM_L_X92Y114_SLICE_X145Y114_AQ),
.I1(CLBLM_R_X93Y119_SLICE_X147Y119_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X92Y114_SLICE_X144Y114_A5Q),
.I4(CLBLM_L_X92Y114_SLICE_X144Y114_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y114_SLICE_X144Y114_CO5),
.O6(CLBLM_L_X92Y114_SLICE_X144Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y114_SLICE_X144Y114_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y113_SLICE_X143Y113_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X144Y114_BO5),
.O6(CLBLM_L_X92Y114_SLICE_X144Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000099990000)
  ) CLBLM_L_X92Y114_SLICE_X144Y114_ALUT (
.I0(CLBLM_L_X92Y114_SLICE_X144Y114_B5Q),
.I1(CLBLM_L_X90Y113_SLICE_X143Y113_A5Q),
.I2(CLBLM_L_X90Y114_SLICE_X143Y114_CO6),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X144Y114_AO5),
.O6(CLBLM_L_X92Y114_SLICE_X144Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y114_SLICE_X145Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y114_SLICE_X145Y114_AO5),
.Q(CLBLM_L_X92Y114_SLICE_X145Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y114_SLICE_X145Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y114_SLICE_X145Y114_AO6),
.Q(CLBLM_L_X92Y114_SLICE_X145Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y114_SLICE_X145Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X145Y114_DO5),
.O6(CLBLM_L_X92Y114_SLICE_X145Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y114_SLICE_X145Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X145Y114_CO5),
.O6(CLBLM_L_X92Y114_SLICE_X145Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y114_SLICE_X145Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X145Y114_BO5),
.O6(CLBLM_L_X92Y114_SLICE_X145Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_L_X92Y114_SLICE_X145Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y114_SLICE_X145Y114_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y113_SLICE_X145Y113_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y114_SLICE_X145Y114_AO5),
.O6(CLBLM_L_X92Y114_SLICE_X145Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y115_SLICE_X144Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y115_SLICE_X144Y115_DO5),
.O6(CLBLM_L_X92Y115_SLICE_X144Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y115_SLICE_X144Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y115_SLICE_X144Y115_CO5),
.O6(CLBLM_L_X92Y115_SLICE_X144Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y115_SLICE_X144Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y115_SLICE_X144Y115_BO5),
.O6(CLBLM_L_X92Y115_SLICE_X144Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y115_SLICE_X144Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y115_SLICE_X144Y115_AO5),
.O6(CLBLM_L_X92Y115_SLICE_X144Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y115_SLICE_X145Y115_AO5),
.Q(CLBLM_L_X92Y115_SLICE_X145Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y115_SLICE_X145Y115_BO5),
.Q(CLBLM_L_X92Y115_SLICE_X145Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y115_SLICE_X145Y115_AO6),
.Q(CLBLM_L_X92Y115_SLICE_X145Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y115_SLICE_X145Y115_BO6),
.Q(CLBLM_L_X92Y115_SLICE_X145Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h73437f4f70407c4c)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_DLUT (
.I0(CLBLM_L_X92Y115_SLICE_X145Y115_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y116_SLICE_X146Y116_CO6),
.I4(CLBLM_L_X94Y116_SLICE_X149Y116_A5Q),
.I5(CLBLM_L_X90Y114_SLICE_X143Y114_DO6),
.O5(CLBLM_L_X92Y115_SLICE_X145Y115_DO5),
.O6(CLBLM_L_X92Y115_SLICE_X145Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3276bafe105498dc)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X90Y114_SLICE_X142Y114_DO6),
.I3(CLBLM_R_X93Y117_SLICE_X146Y117_A5Q),
.I4(CLBLM_L_X92Y115_SLICE_X145Y115_AQ),
.I5(CLBLM_R_X93Y117_SLICE_X146Y117_CO6),
.O5(CLBLM_L_X92Y115_SLICE_X145Y115_CO5),
.O6(CLBLM_L_X92Y115_SLICE_X145Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500cc003300)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_BLUT (
.I0(CLBLM_L_X92Y115_SLICE_X145Y115_DO6),
.I1(CLBLM_R_X93Y115_SLICE_X147Y115_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y114_SLICE_X143Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y115_SLICE_X145Y115_BO5),
.O6(CLBLM_L_X92Y115_SLICE_X145Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_L_X92Y115_SLICE_X145Y115_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y114_SLICE_X149Y114_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y115_SLICE_X145Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y115_SLICE_X145Y115_AO5),
.O6(CLBLM_L_X92Y115_SLICE_X145Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X144Y116_AO5),
.Q(CLBLM_L_X92Y116_SLICE_X144Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X144Y116_BO5),
.Q(CLBLM_L_X92Y116_SLICE_X144Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X144Y116_AO6),
.Q(CLBLM_L_X92Y116_SLICE_X144Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X144Y116_BO6),
.Q(CLBLM_L_X92Y116_SLICE_X144Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X92Y116_SLICE_X144Y116_AQ),
.I2(CLBLM_L_X92Y116_SLICE_X144Y116_BQ),
.I3(CLBLM_L_X92Y119_SLICE_X144Y119_CQ),
.I4(CLBLM_L_X92Y116_SLICE_X144Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y116_SLICE_X144Y116_DO5),
.O6(CLBLM_L_X92Y116_SLICE_X144Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h330f330fffaa00aa)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_CLUT (
.I0(CLBLM_R_X93Y120_SLICE_X146Y120_DO6),
.I1(CLBLM_L_X90Y116_SLICE_X143Y116_AQ),
.I2(CLBLM_L_X90Y116_SLICE_X143Y116_C5Q),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X92Y116_SLICE_X144Y116_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y116_SLICE_X144Y116_CO5),
.O6(CLBLM_L_X92Y116_SLICE_X144Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y116_SLICE_X144Y116_AQ),
.I3(1'b1),
.I4(CLBLM_L_X92Y116_SLICE_X144Y116_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y116_SLICE_X144Y116_BO5),
.O6(CLBLM_L_X92Y116_SLICE_X144Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_L_X92Y116_SLICE_X144Y116_ALUT (
.I0(CLBLM_L_X90Y118_SLICE_X142Y118_B5Q),
.I1(CLBLM_L_X92Y119_SLICE_X144Y119_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y116_SLICE_X144Y116_AO5),
.O6(CLBLM_L_X92Y116_SLICE_X144Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X145Y116_AO5),
.Q(CLBLM_L_X92Y116_SLICE_X145Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X145Y116_BO5),
.Q(CLBLM_L_X92Y116_SLICE_X145Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X145Y116_AO6),
.Q(CLBLM_L_X92Y116_SLICE_X145Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y116_SLICE_X145Y116_BO6),
.Q(CLBLM_L_X92Y116_SLICE_X145Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_DLUT (
.I0(CLBLM_L_X90Y116_SLICE_X142Y116_AQ),
.I1(CLBLM_L_X90Y116_SLICE_X142Y116_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X92Y116_SLICE_X145Y116_BQ),
.I4(CLBLM_L_X92Y116_SLICE_X145Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y116_SLICE_X145Y116_DO5),
.O6(CLBLM_L_X92Y116_SLICE_X145Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h737f434f707c404c)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_CLUT (
.I0(CLBLM_L_X90Y115_SLICE_X143Y115_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X92Y116_SLICE_X145Y116_A5Q),
.I4(CLBLM_L_X92Y116_SLICE_X145Y116_DO6),
.I5(CLBLM_L_X90Y118_SLICE_X142Y118_DO6),
.O5(CLBLM_L_X92Y116_SLICE_X145Y116_CO5),
.O6(CLBLM_L_X92Y116_SLICE_X145Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_BLUT (
.I0(CLBLM_L_X90Y116_SLICE_X142Y116_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y116_SLICE_X145Y116_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y116_SLICE_X145Y116_BO5),
.O6(CLBLM_L_X92Y116_SLICE_X145Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0099009900)
  ) CLBLM_L_X92Y116_SLICE_X145Y116_ALUT (
.I0(CLBLM_L_X92Y116_SLICE_X145Y116_B5Q),
.I1(CLBLM_R_X89Y115_SLICE_X141Y115_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X100Y116_SLICE_X157Y116_CO6),
.I5(1'b1),
.O5(CLBLM_L_X92Y116_SLICE_X145Y116_AO5),
.O6(CLBLM_L_X92Y116_SLICE_X145Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y118_SLICE_X144Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y118_SLICE_X144Y118_AO5),
.Q(CLBLM_L_X92Y118_SLICE_X144Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y118_SLICE_X144Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y118_SLICE_X144Y118_AO6),
.Q(CLBLM_L_X92Y118_SLICE_X144Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y118_SLICE_X144Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X144Y118_DO5),
.O6(CLBLM_L_X92Y118_SLICE_X144Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y118_SLICE_X144Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X144Y118_CO5),
.O6(CLBLM_L_X92Y118_SLICE_X144Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeeb1441ebbe4114)
  ) CLBLM_L_X92Y118_SLICE_X144Y118_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X89Y118_SLICE_X141Y118_A5Q),
.I2(CLBLM_R_X89Y115_SLICE_X141Y115_BQ),
.I3(CLBLM_R_X89Y118_SLICE_X141Y118_AQ),
.I4(CLBLM_R_X97Y119_SLICE_X152Y119_CQ),
.I5(CLBLM_L_X92Y118_SLICE_X144Y118_A5Q),
.O5(CLBLM_L_X92Y118_SLICE_X144Y118_BO5),
.O6(CLBLM_L_X92Y118_SLICE_X144Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_L_X92Y118_SLICE_X144Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X89Y115_SLICE_X141Y115_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y119_SLICE_X144Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X144Y118_AO5),
.O6(CLBLM_L_X92Y118_SLICE_X144Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y118_SLICE_X145Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X145Y118_DO5),
.O6(CLBLM_L_X92Y118_SLICE_X145Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y118_SLICE_X145Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X145Y118_CO5),
.O6(CLBLM_L_X92Y118_SLICE_X145Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y118_SLICE_X145Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X145Y118_BO5),
.O6(CLBLM_L_X92Y118_SLICE_X145Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y118_SLICE_X145Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y118_SLICE_X145Y118_AO5),
.O6(CLBLM_L_X92Y118_SLICE_X145Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X144Y119_BO5),
.Q(CLBLM_L_X92Y119_SLICE_X144Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X144Y119_CO5),
.Q(CLBLM_L_X92Y119_SLICE_X144Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X144Y119_AO6),
.Q(CLBLM_L_X92Y119_SLICE_X144Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X144Y119_CO6),
.Q(CLBLM_L_X92Y119_SLICE_X144Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y119_SLICE_X144Y119_DO5),
.O6(CLBLM_L_X92Y119_SLICE_X144Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300f0000f00)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y116_SLICE_X144Y116_CO6),
.I2(CLBLM_L_X92Y119_SLICE_X145Y119_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y120_SLICE_X143Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y119_SLICE_X144Y119_CO5),
.O6(CLBLM_L_X92Y119_SLICE_X144Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acc00cc00)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_BLUT (
.I0(CLBLM_L_X92Y118_SLICE_X144Y118_AQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y119_SLICE_X144Y119_AQ),
.I3(CLBLM_L_X92Y120_SLICE_X145Y120_C5Q),
.I4(CLBLM_L_X92Y119_SLICE_X144Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y119_SLICE_X144Y119_BO5),
.O6(CLBLM_L_X92Y119_SLICE_X144Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb00c80073004000)
  ) CLBLM_L_X92Y119_SLICE_X144Y119_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X92Y119_SLICE_X144Y119_BO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y123_SLICE_X143Y123_DO6),
.I5(CLBLM_L_X92Y121_SLICE_X144Y121_A5Q),
.O5(CLBLM_L_X92Y119_SLICE_X144Y119_AO5),
.O6(CLBLM_L_X92Y119_SLICE_X144Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X145Y119_AO5),
.Q(CLBLM_L_X92Y119_SLICE_X145Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X145Y119_BO5),
.Q(CLBLM_L_X92Y119_SLICE_X145Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X145Y119_AO6),
.Q(CLBLM_L_X92Y119_SLICE_X145Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y119_SLICE_X145Y119_BO6),
.Q(CLBLM_L_X92Y119_SLICE_X145Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_DLUT (
.I0(CLBLM_R_X93Y124_SLICE_X147Y124_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(1'b1),
.I3(CLBLM_L_X92Y119_SLICE_X145Y119_BQ),
.I4(CLBLM_L_X92Y119_SLICE_X145Y119_B5Q),
.I5(CLBLM_L_X90Y119_SLICE_X143Y119_BQ),
.O5(CLBLM_L_X92Y119_SLICE_X145Y119_DO5),
.O6(CLBLM_L_X92Y119_SLICE_X145Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_CLUT (
.I0(CLBLM_L_X92Y118_SLICE_X144Y118_AQ),
.I1(CLBLM_L_X92Y120_SLICE_X145Y120_C5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y120_SLICE_X153Y120_C5Q),
.I4(CLBLM_L_X92Y119_SLICE_X144Y119_AQ),
.I5(CLBLM_L_X92Y119_SLICE_X144Y119_A5Q),
.O5(CLBLM_L_X92Y119_SLICE_X145Y119_CO5),
.O6(CLBLM_L_X92Y119_SLICE_X145Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_L_X90Y119_SLICE_X143Y119_BQ),
.I4(CLBLM_L_X92Y119_SLICE_X145Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y119_SLICE_X145Y119_BO5),
.O6(CLBLM_L_X92Y119_SLICE_X145Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc000f000f00)
  ) CLBLM_L_X92Y119_SLICE_X145Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y119_SLICE_X145Y119_A5Q),
.I2(CLBLM_L_X92Y115_SLICE_X145Y115_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y119_SLICE_X145Y119_AO5),
.O6(CLBLM_L_X92Y119_SLICE_X145Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X144Y120_AO5),
.Q(CLBLM_L_X92Y120_SLICE_X144Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X144Y120_BO5),
.Q(CLBLM_L_X92Y120_SLICE_X144Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X144Y120_AO6),
.Q(CLBLM_L_X92Y120_SLICE_X144Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X144Y120_BO6),
.Q(CLBLM_L_X92Y120_SLICE_X144Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_DLUT (
.I0(CLBLM_L_X92Y120_SLICE_X144Y120_BQ),
.I1(1'b1),
.I2(CLBLM_R_X93Y120_SLICE_X146Y120_AQ),
.I3(CLBLM_L_X90Y122_SLICE_X143Y122_C5Q),
.I4(CLBLM_L_X92Y120_SLICE_X144Y120_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y120_SLICE_X144Y120_DO5),
.O6(CLBLM_L_X92Y120_SLICE_X144Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bb11bbfafa5050)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X90Y120_SLICE_X143Y120_A5Q),
.I2(CLBLM_R_X93Y124_SLICE_X147Y124_DO6),
.I3(CLBLM_L_X92Y120_SLICE_X144Y120_A5Q),
.I4(CLBLM_L_X92Y120_SLICE_X144Y120_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y120_SLICE_X144Y120_CO5),
.O6(CLBLM_L_X92Y120_SLICE_X144Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_BLUT (
.I0(CLBLM_R_X93Y120_SLICE_X146Y120_AQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y120_SLICE_X144Y120_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y120_SLICE_X144Y120_BO5),
.O6(CLBLM_L_X92Y120_SLICE_X144Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_L_X92Y120_SLICE_X144Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y120_SLICE_X144Y120_A5Q),
.I2(CLBLM_L_X90Y120_SLICE_X142Y120_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y120_SLICE_X144Y120_AO5),
.O6(CLBLM_L_X92Y120_SLICE_X144Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X145Y120_BO5),
.Q(CLBLM_L_X92Y120_SLICE_X145Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X145Y120_CO5),
.Q(CLBLM_L_X92Y120_SLICE_X145Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X145Y120_AO6),
.Q(CLBLM_L_X92Y120_SLICE_X145Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y120_SLICE_X145Y120_CO6),
.Q(CLBLM_L_X92Y120_SLICE_X145Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_DLUT (
.I0(CLBLM_R_X97Y120_SLICE_X153Y120_CQ),
.I1(CLBLM_L_X92Y120_SLICE_X145Y120_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y120_SLICE_X145Y120_A5Q),
.I4(CLBLM_L_X92Y120_SLICE_X145Y120_AQ),
.I5(CLBLM_L_X94Y121_SLICE_X148Y121_C5Q),
.O5(CLBLM_L_X92Y120_SLICE_X145Y120_DO5),
.O6(CLBLM_L_X92Y120_SLICE_X145Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X92Y118_SLICE_X144Y118_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y120_SLICE_X145Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y120_SLICE_X145Y120_CO5),
.O6(CLBLM_L_X92Y120_SLICE_X145Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acc00cc00)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_BLUT (
.I0(CLBLM_L_X92Y120_SLICE_X145Y120_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y120_SLICE_X145Y120_AQ),
.I3(CLBLM_L_X94Y121_SLICE_X148Y121_C5Q),
.I4(CLBLM_L_X92Y120_SLICE_X145Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y120_SLICE_X145Y120_BO5),
.O6(CLBLM_L_X92Y120_SLICE_X145Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heee22e2200000000)
  ) CLBLM_L_X92Y120_SLICE_X145Y120_ALUT (
.I0(CLBLM_L_X92Y121_SLICE_X145Y121_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y120_SLICE_X145Y120_BO6),
.I4(CLBLM_L_X92Y119_SLICE_X145Y119_A5Q),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X92Y120_SLICE_X145Y120_AO5),
.O6(CLBLM_L_X92Y120_SLICE_X145Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X144Y121_AO5),
.Q(CLBLM_L_X92Y121_SLICE_X144Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X144Y121_DO5),
.Q(CLBLM_L_X92Y121_SLICE_X144Y121_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X144Y121_AO6),
.Q(CLBLM_L_X92Y121_SLICE_X144Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X144Y121_BO6),
.Q(CLBLM_L_X92Y121_SLICE_X144Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X144Y121_CO6),
.Q(CLBLM_L_X92Y121_SLICE_X144Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X144Y121_DO6),
.Q(CLBLM_L_X92Y121_SLICE_X144Y121_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc030c03050a0a050)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_DLUT (
.I0(CLBLM_L_X92Y119_SLICE_X144Y119_A5Q),
.I1(CLBLM_L_X92Y120_SLICE_X145Y120_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y117_SLICE_X146Y117_A5Q),
.I4(CLBLM_L_X92Y122_SLICE_X145Y122_CQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y121_SLICE_X144Y121_DO5),
.O6(CLBLM_L_X92Y121_SLICE_X144Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5dda08800000000)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X92Y121_SLICE_X145Y121_AO6),
.I2(CLBLM_L_X90Y114_SLICE_X142Y114_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X90Y125_SLICE_X142Y125_BO6),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X92Y121_SLICE_X144Y121_CO5),
.O6(CLBLM_L_X92Y121_SLICE_X144Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0cc00088888888)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_BLUT (
.I0(CLBLM_L_X92Y122_SLICE_X144Y122_DO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y121_SLICE_X146Y121_AQ),
.I4(CLBLM_R_X93Y121_SLICE_X146Y121_BO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y121_SLICE_X144Y121_BO5),
.O6(CLBLM_L_X92Y121_SLICE_X144Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_L_X92Y121_SLICE_X144Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y121_SLICE_X144Y121_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y121_SLICE_X146Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y121_SLICE_X144Y121_AO5),
.O6(CLBLM_L_X92Y121_SLICE_X144Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X145Y121_BO5),
.Q(CLBLM_L_X92Y121_SLICE_X145Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X145Y121_CO5),
.Q(CLBLM_L_X92Y121_SLICE_X145Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X145Y121_AO5),
.Q(CLBLM_L_X92Y121_SLICE_X145Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X145Y121_BO6),
.Q(CLBLM_L_X92Y121_SLICE_X145Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y121_SLICE_X145Y121_CO6),
.Q(CLBLM_L_X92Y121_SLICE_X145Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_DLUT (
.I0(CLBLM_L_X92Y121_SLICE_X144Y121_CQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X92Y121_SLICE_X145Y121_BQ),
.I3(CLBLM_L_X92Y121_SLICE_X145Y121_AQ),
.I4(CLBLM_L_X92Y121_SLICE_X145Y121_B5Q),
.I5(CLBLM_L_X92Y121_SLICE_X144Y121_DQ),
.O5(CLBLM_L_X92Y121_SLICE_X145Y121_DO5),
.O6(CLBLM_L_X92Y121_SLICE_X145Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa005500c300c300)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_CLUT (
.I0(CLBLM_L_X92Y121_SLICE_X144Y121_DQ),
.I1(CLBLM_L_X92Y121_SLICE_X145Y121_CQ),
.I2(CLBLM_R_X93Y121_SLICE_X147Y121_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y121_SLICE_X148Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y121_SLICE_X145Y121_CO5),
.O6(CLBLM_L_X92Y121_SLICE_X145Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_BLUT (
.I0(CLBLM_L_X92Y121_SLICE_X145Y121_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y121_SLICE_X144Y121_CQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y121_SLICE_X145Y121_BO5),
.O6(CLBLM_L_X92Y121_SLICE_X145Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_L_X92Y121_SLICE_X145Y121_ALUT (
.I0(CLBLM_L_X92Y121_SLICE_X145Y121_B5Q),
.I1(CLBLM_L_X92Y121_SLICE_X145Y121_BQ),
.I2(CLBLM_L_X92Y121_SLICE_X145Y121_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y121_SLICE_X144Y121_CQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y121_SLICE_X145Y121_AO5),
.O6(CLBLM_L_X92Y121_SLICE_X145Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X144Y122_BO5),
.Q(CLBLM_L_X92Y122_SLICE_X144Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X144Y122_CO5),
.Q(CLBLM_L_X92Y122_SLICE_X144Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X144Y122_AO5),
.Q(CLBLM_L_X92Y122_SLICE_X144Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X144Y122_BO6),
.Q(CLBLM_L_X92Y122_SLICE_X144Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X144Y122_CO6),
.Q(CLBLM_L_X92Y122_SLICE_X144Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12ed21ed21de12)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_DLUT (
.I0(CLBLM_L_X92Y122_SLICE_X144Y122_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X92Y122_SLICE_X144Y122_AQ),
.I3(CLBLM_L_X92Y122_SLICE_X145Y122_CQ),
.I4(CLBLM_L_X92Y122_SLICE_X144Y122_B5Q),
.I5(CLBLM_L_X90Y122_SLICE_X142Y122_BQ),
.O5(CLBLM_L_X92Y122_SLICE_X144Y122_DO5),
.O6(CLBLM_L_X92Y122_SLICE_X144Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha500a500cc003300)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_CLUT (
.I0(CLBLM_L_X90Y124_SLICE_X143Y124_C5Q),
.I1(CLBLM_L_X92Y122_SLICE_X144Y122_CQ),
.I2(CLBLM_L_X90Y120_SLICE_X142Y120_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X90Y119_SLICE_X143Y119_CQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X144Y122_CO5),
.O6(CLBLM_L_X92Y122_SLICE_X144Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y122_SLICE_X144Y122_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y122_SLICE_X142Y122_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X144Y122_BO5),
.O6(CLBLM_L_X92Y122_SLICE_X144Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_L_X92Y122_SLICE_X144Y122_ALUT (
.I0(CLBLM_L_X92Y122_SLICE_X144Y122_B5Q),
.I1(CLBLM_L_X90Y122_SLICE_X142Y122_BQ),
.I2(CLBLM_L_X92Y122_SLICE_X144Y122_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y122_SLICE_X144Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X144Y122_AO5),
.O6(CLBLM_L_X92Y122_SLICE_X144Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X145Y122_BO5),
.Q(CLBLM_L_X92Y122_SLICE_X145Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X145Y122_CO5),
.Q(CLBLM_L_X92Y122_SLICE_X145Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X145Y122_AO5),
.Q(CLBLM_L_X92Y122_SLICE_X145Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X145Y122_BO6),
.Q(CLBLM_L_X92Y122_SLICE_X145Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y122_SLICE_X145Y122_CO6),
.Q(CLBLM_L_X92Y122_SLICE_X145Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X145Y122_DO5),
.O6(CLBLM_L_X92Y122_SLICE_X145Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88448844c0c00c0c)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_CLUT (
.I0(CLBLM_R_X93Y121_SLICE_X146Y121_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y122_SLICE_X147Y122_A5Q),
.I3(CLBLM_L_X92Y121_SLICE_X145Y121_C5Q),
.I4(CLBLM_L_X92Y121_SLICE_X144Y121_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X145Y122_CO5),
.O6(CLBLM_L_X92Y122_SLICE_X145Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cc00cc00)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y120_SLICE_X140Y120_AQ),
.I3(CLBLM_R_X93Y122_SLICE_X146Y122_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X145Y122_BO5),
.O6(CLBLM_L_X92Y122_SLICE_X145Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996aaaa0000)
  ) CLBLM_L_X92Y122_SLICE_X145Y122_ALUT (
.I0(CLBLM_L_X92Y122_SLICE_X145Y122_B5Q),
.I1(CLBLM_R_X93Y122_SLICE_X146Y122_AQ),
.I2(CLBLM_L_X92Y122_SLICE_X145Y122_AQ),
.I3(CLBLM_L_X92Y123_SLICE_X145Y123_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X92Y122_SLICE_X145Y122_AO5),
.O6(CLBLM_L_X92Y122_SLICE_X145Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X144Y123_AO5),
.Q(CLBLM_L_X92Y123_SLICE_X144Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X144Y123_DO5),
.Q(CLBLM_L_X92Y123_SLICE_X144Y123_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X144Y123_AO6),
.Q(CLBLM_L_X92Y123_SLICE_X144Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X144Y123_BO6),
.Q(CLBLM_L_X92Y123_SLICE_X144Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X144Y123_CO6),
.Q(CLBLM_L_X92Y123_SLICE_X144Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X144Y123_DO6),
.Q(CLBLM_L_X92Y123_SLICE_X144Y123_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00a0a88228822)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y123_SLICE_X144Y123_DQ),
.I2(CLBLM_L_X92Y123_SLICE_X145Y123_B5Q),
.I3(CLBLM_L_X92Y122_SLICE_X145Y122_AQ),
.I4(CLBLM_L_X92Y124_SLICE_X145Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y123_SLICE_X144Y123_DO5),
.O6(CLBLM_L_X92Y123_SLICE_X144Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha808a808aaaa0000)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y123_SLICE_X147Y123_AO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y123_SLICE_X144Y123_A5Q),
.I4(CLBLM_L_X92Y124_SLICE_X144Y124_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y123_SLICE_X144Y123_CO5),
.O6(CLBLM_L_X92Y123_SLICE_X144Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000c0c0a0a0a0a0)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_BLUT (
.I0(CLBLM_L_X90Y126_SLICE_X143Y126_DO6),
.I1(CLBLM_R_X93Y123_SLICE_X146Y123_AO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y123_SLICE_X144Y123_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y123_SLICE_X144Y123_BO5),
.O6(CLBLM_L_X92Y123_SLICE_X144Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X92Y123_SLICE_X144Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y123_SLICE_X144Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X92Y121_SLICE_X144Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y123_SLICE_X144Y123_AO5),
.O6(CLBLM_L_X92Y123_SLICE_X144Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X145Y123_AO5),
.Q(CLBLM_L_X92Y123_SLICE_X145Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X145Y123_DO5),
.Q(CLBLM_L_X92Y123_SLICE_X145Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X145Y123_AO6),
.Q(CLBLM_L_X92Y123_SLICE_X145Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X145Y123_BO6),
.Q(CLBLM_L_X92Y123_SLICE_X145Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y123_SLICE_X145Y123_CO6),
.Q(CLBLM_L_X92Y123_SLICE_X145Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33ca0a0a0a0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y123_SLICE_X145Y123_CQ),
.I2(CLBLM_R_X93Y122_SLICE_X146Y122_A5Q),
.I3(CLBLM_R_X93Y123_SLICE_X146Y123_BQ),
.I4(CLBLM_L_X92Y123_SLICE_X145Y123_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y123_SLICE_X145Y123_DO5),
.O6(CLBLM_L_X92Y123_SLICE_X145Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa228800a0a0a0a0)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X90Y126_SLICE_X142Y126_DO6),
.I3(CLBLM_L_X92Y123_SLICE_X145Y123_A5Q),
.I4(CLBLM_L_X92Y123_SLICE_X145Y123_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y123_SLICE_X145Y123_CO5),
.O6(CLBLM_L_X92Y123_SLICE_X145Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf070b030c0408000)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y123_SLICE_X145Y123_AQ),
.I4(CLBLM_L_X92Y122_SLICE_X145Y122_AO6),
.I5(CLBLM_R_X89Y123_SLICE_X140Y123_DO6),
.O5(CLBLM_L_X92Y123_SLICE_X145Y123_BO5),
.O6(CLBLM_L_X92Y123_SLICE_X145Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X92Y123_SLICE_X145Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X92Y123_SLICE_X145Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X92Y123_SLICE_X144Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y123_SLICE_X145Y123_AO5),
.O6(CLBLM_L_X92Y123_SLICE_X145Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y124_SLICE_X144Y124_BO5),
.Q(CLBLM_L_X92Y124_SLICE_X144Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y124_SLICE_X144Y124_CO5),
.Q(CLBLM_L_X92Y124_SLICE_X144Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y124_SLICE_X144Y124_AO6),
.Q(CLBLM_L_X92Y124_SLICE_X144Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y124_SLICE_X144Y124_CO6),
.Q(CLBLM_L_X92Y124_SLICE_X144Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5aa5cccca55a)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_DLUT (
.I0(CLBLM_L_X92Y124_SLICE_X144Y124_C5Q),
.I1(CLBLM_L_X92Y124_SLICE_X145Y124_AQ),
.I2(CLBLM_L_X92Y124_SLICE_X144Y124_AQ),
.I3(CLBLM_L_X92Y124_SLICE_X144Y124_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X92Y124_SLICE_X144Y124_CQ),
.O5(CLBLM_L_X92Y124_SLICE_X144Y124_DO5),
.O6(CLBLM_L_X92Y124_SLICE_X144Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y124_SLICE_X144Y124_CQ),
.I2(CLBLM_L_X92Y124_SLICE_X144Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y124_SLICE_X144Y124_CO5),
.O6(CLBLM_L_X92Y124_SLICE_X144Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_BLUT (
.I0(CLBLM_L_X92Y124_SLICE_X144Y124_AQ),
.I1(CLBLM_L_X92Y124_SLICE_X144Y124_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y124_SLICE_X144Y124_CQ),
.I4(CLBLM_L_X92Y124_SLICE_X144Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y124_SLICE_X144Y124_BO5),
.O6(CLBLM_L_X92Y124_SLICE_X144Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e02020e020e020)
  ) CLBLM_L_X92Y124_SLICE_X144Y124_ALUT (
.I0(CLBLM_L_X90Y130_SLICE_X142Y130_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y124_SLICE_X144Y124_BO6),
.I4(CLBLM_L_X90Y123_SLICE_X142Y123_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y124_SLICE_X144Y124_AO5),
.O6(CLBLM_L_X92Y124_SLICE_X144Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y124_SLICE_X145Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y124_SLICE_X145Y124_AO5),
.Q(CLBLM_L_X92Y124_SLICE_X145Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y124_SLICE_X145Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y124_SLICE_X145Y124_AO6),
.Q(CLBLM_L_X92Y124_SLICE_X145Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y124_SLICE_X145Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y124_SLICE_X145Y124_DO5),
.O6(CLBLM_L_X92Y124_SLICE_X145Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y124_SLICE_X145Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y124_SLICE_X145Y124_CO5),
.O6(CLBLM_L_X92Y124_SLICE_X145Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y124_SLICE_X145Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y124_SLICE_X145Y124_BO5),
.O6(CLBLM_L_X92Y124_SLICE_X145Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05050c030c030)
  ) CLBLM_L_X92Y124_SLICE_X145Y124_ALUT (
.I0(CLBLM_R_X93Y123_SLICE_X146Y123_CQ),
.I1(CLBLM_R_X93Y123_SLICE_X146Y123_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y124_SLICE_X145Y124_AQ),
.I4(CLBLM_L_X92Y122_SLICE_X145Y122_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y124_SLICE_X145Y124_AO5),
.O6(CLBLM_L_X92Y124_SLICE_X145Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_DO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_CO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_BO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y125_SLICE_X144Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X144Y125_AO5),
.O6(CLBLM_L_X92Y125_SLICE_X144Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y125_SLICE_X145Y125_BO5),
.Q(CLBLM_L_X92Y125_SLICE_X145Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y125_SLICE_X145Y125_CO5),
.Q(CLBLM_L_X92Y125_SLICE_X145Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y125_SLICE_X145Y125_AO6),
.Q(CLBLM_L_X92Y125_SLICE_X145Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y125_SLICE_X145Y125_CO6),
.Q(CLBLM_L_X92Y125_SLICE_X145Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_DLUT (
.I0(CLBLM_L_X92Y125_SLICE_X145Y125_C5Q),
.I1(CLBLM_L_X92Y125_SLICE_X145Y125_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y125_SLICE_X145Y125_A5Q),
.I4(CLBLM_L_X92Y125_SLICE_X145Y125_AQ),
.I5(CLBLM_L_X90Y124_SLICE_X143Y124_CQ),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_DO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y125_SLICE_X145Y125_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y125_SLICE_X145Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_CO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_BLUT (
.I0(CLBLM_L_X92Y125_SLICE_X145Y125_AQ),
.I1(CLBLM_L_X92Y125_SLICE_X145Y125_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y125_SLICE_X145Y125_CQ),
.I4(CLBLM_L_X92Y125_SLICE_X145Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_BO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a05000c0c0c0c0)
  ) CLBLM_L_X92Y125_SLICE_X145Y125_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X94Y126_SLICE_X149Y126_AO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y125_SLICE_X145Y125_BO6),
.I4(CLBLM_R_X93Y127_SLICE_X146Y127_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y125_SLICE_X145Y125_AO5),
.O6(CLBLM_L_X92Y125_SLICE_X145Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y126_SLICE_X144Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y126_SLICE_X145Y126_AO5),
.Q(CLBLM_L_X92Y126_SLICE_X144Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y126_SLICE_X144Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X144Y126_DO5),
.O6(CLBLM_L_X92Y126_SLICE_X144Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y126_SLICE_X144Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X144Y126_CO5),
.O6(CLBLM_L_X92Y126_SLICE_X144Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y126_SLICE_X144Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X144Y126_BO5),
.O6(CLBLM_L_X92Y126_SLICE_X144Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y126_SLICE_X144Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X144Y126_AO5),
.O6(CLBLM_L_X92Y126_SLICE_X144Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y126_SLICE_X145Y126_BO5),
.Q(CLBLM_L_X92Y126_SLICE_X145Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y126_SLICE_X145Y126_CO5),
.Q(CLBLM_L_X92Y126_SLICE_X145Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y126_SLICE_X145Y126_BO6),
.Q(CLBLM_L_X92Y126_SLICE_X145Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y126_SLICE_X145Y126_CO6),
.Q(CLBLM_L_X92Y126_SLICE_X145Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_DLUT (
.I0(CLBLM_L_X92Y126_SLICE_X144Y126_AQ),
.I1(CLBLM_L_X92Y126_SLICE_X145Y126_CQ),
.I2(CLBLM_L_X92Y126_SLICE_X145Y126_BQ),
.I3(CLBLM_R_X93Y127_SLICE_X146Y127_CQ),
.I4(CLBLM_L_X92Y126_SLICE_X145Y126_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y126_SLICE_X145Y126_DO5),
.O6(CLBLM_L_X92Y126_SLICE_X145Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha050a050c0c03030)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_CLUT (
.I0(CLBLM_L_X90Y125_SLICE_X143Y125_BQ),
.I1(CLBLM_L_X92Y126_SLICE_X145Y126_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y125_SLICE_X141Y125_A5Q),
.I4(CLBLM_R_X89Y126_SLICE_X141Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X145Y126_CO5),
.O6(CLBLM_L_X92Y126_SLICE_X145Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y126_SLICE_X145Y126_BQ),
.I2(1'b1),
.I3(CLBLM_R_X93Y127_SLICE_X146Y127_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X145Y126_BO5),
.O6(CLBLM_L_X92Y126_SLICE_X145Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_L_X92Y126_SLICE_X145Y126_ALUT (
.I0(CLBLM_L_X92Y126_SLICE_X145Y126_B5Q),
.I1(CLBLM_L_X92Y126_SLICE_X145Y126_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y127_SLICE_X146Y127_CQ),
.I4(CLBLM_L_X92Y126_SLICE_X144Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y126_SLICE_X145Y126_AO5),
.O6(CLBLM_L_X92Y126_SLICE_X145Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y127_SLICE_X144Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X144Y127_DO5),
.O6(CLBLM_L_X92Y127_SLICE_X144Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y127_SLICE_X144Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X144Y127_CO5),
.O6(CLBLM_L_X92Y127_SLICE_X144Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y127_SLICE_X144Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X144Y127_BO5),
.O6(CLBLM_L_X92Y127_SLICE_X144Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y127_SLICE_X144Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X144Y127_AO5),
.O6(CLBLM_L_X92Y127_SLICE_X144Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y127_SLICE_X145Y127_BO5),
.Q(CLBLM_L_X92Y127_SLICE_X145Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y127_SLICE_X145Y127_AO5),
.Q(CLBLM_L_X92Y127_SLICE_X145Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y127_SLICE_X145Y127_BO6),
.Q(CLBLM_L_X92Y127_SLICE_X145Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X145Y127_DO5),
.O6(CLBLM_L_X92Y127_SLICE_X145Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_CLUT (
.I0(CLBLM_R_X93Y127_SLICE_X146Y127_BQ),
.I1(CLBLM_L_X90Y125_SLICE_X143Y125_CQ),
.I2(CLBLM_L_X92Y127_SLICE_X145Y127_BQ),
.I3(CLBLM_L_X92Y127_SLICE_X145Y127_AQ),
.I4(CLBLM_L_X92Y127_SLICE_X145Y127_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y127_SLICE_X145Y127_CO5),
.O6(CLBLM_L_X92Y127_SLICE_X145Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_BLUT (
.I0(CLBLM_L_X92Y127_SLICE_X145Y127_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y127_SLICE_X146Y127_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X145Y127_BO5),
.O6(CLBLM_L_X92Y127_SLICE_X145Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acc00cc00)
  ) CLBLM_L_X92Y127_SLICE_X145Y127_ALUT (
.I0(CLBLM_L_X92Y127_SLICE_X145Y127_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y127_SLICE_X145Y127_AQ),
.I3(CLBLM_L_X92Y127_SLICE_X145Y127_B5Q),
.I4(CLBLM_R_X93Y127_SLICE_X146Y127_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y127_SLICE_X145Y127_AO5),
.O6(CLBLM_L_X92Y127_SLICE_X145Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y128_SLICE_X144Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y128_SLICE_X144Y128_DO5),
.O6(CLBLM_L_X92Y128_SLICE_X144Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y128_SLICE_X144Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y128_SLICE_X144Y128_CO5),
.O6(CLBLM_L_X92Y128_SLICE_X144Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y128_SLICE_X144Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y128_SLICE_X144Y128_BO5),
.O6(CLBLM_L_X92Y128_SLICE_X144Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y128_SLICE_X144Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y128_SLICE_X144Y128_AO5),
.O6(CLBLM_L_X92Y128_SLICE_X144Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y128_SLICE_X145Y128_BO5),
.Q(CLBLM_L_X92Y128_SLICE_X145Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y128_SLICE_X145Y128_CO5),
.Q(CLBLM_L_X92Y128_SLICE_X145Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y128_SLICE_X145Y128_AO6),
.Q(CLBLM_L_X92Y128_SLICE_X145Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y128_SLICE_X145Y128_CO6),
.Q(CLBLM_L_X92Y128_SLICE_X145Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5aa5a55a)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_DLUT (
.I0(CLBLM_L_X92Y128_SLICE_X145Y128_C5Q),
.I1(CLBLM_L_X90Y125_SLICE_X143Y125_B5Q),
.I2(CLBLM_L_X92Y128_SLICE_X145Y128_CQ),
.I3(CLBLM_L_X92Y128_SLICE_X145Y128_A5Q),
.I4(CLBLM_L_X92Y128_SLICE_X145Y128_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y128_SLICE_X145Y128_DO5),
.O6(CLBLM_L_X92Y128_SLICE_X145Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y128_SLICE_X145Y128_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y128_SLICE_X145Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y128_SLICE_X145Y128_CO5),
.O6(CLBLM_L_X92Y128_SLICE_X145Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996cccc0000)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_BLUT (
.I0(CLBLM_L_X92Y128_SLICE_X145Y128_AQ),
.I1(CLBLM_L_X92Y128_SLICE_X145Y128_C5Q),
.I2(CLBLM_L_X92Y128_SLICE_X145Y128_A5Q),
.I3(CLBLM_L_X92Y128_SLICE_X145Y128_CQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X92Y128_SLICE_X145Y128_BO5),
.O6(CLBLM_L_X92Y128_SLICE_X145Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa005000cc00cc00)
  ) CLBLM_L_X92Y128_SLICE_X145Y128_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X94Y129_SLICE_X148Y129_CO6),
.I2(CLBLM_L_X92Y128_SLICE_X145Y128_BO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y129_SLICE_X146Y129_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X92Y128_SLICE_X145Y128_AO5),
.O6(CLBLM_L_X92Y128_SLICE_X145Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y129_SLICE_X144Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y129_SLICE_X144Y129_DO5),
.O6(CLBLM_L_X92Y129_SLICE_X144Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y129_SLICE_X144Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y129_SLICE_X144Y129_CO5),
.O6(CLBLM_L_X92Y129_SLICE_X144Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y129_SLICE_X144Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y129_SLICE_X144Y129_BO5),
.O6(CLBLM_L_X92Y129_SLICE_X144Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y129_SLICE_X144Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y129_SLICE_X144Y129_AO5),
.O6(CLBLM_L_X92Y129_SLICE_X144Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y129_SLICE_X145Y129_BO5),
.Q(CLBLM_L_X92Y129_SLICE_X145Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y129_SLICE_X145Y129_CO5),
.Q(CLBLM_L_X92Y129_SLICE_X145Y129_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y129_SLICE_X145Y129_AO6),
.Q(CLBLM_L_X92Y129_SLICE_X145Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y129_SLICE_X145Y129_CO6),
.Q(CLBLM_L_X92Y129_SLICE_X145Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_DLUT (
.I0(CLBLM_L_X92Y129_SLICE_X145Y129_C5Q),
.I1(CLBLM_L_X92Y129_SLICE_X145Y129_CQ),
.I2(CLBLM_L_X90Y128_SLICE_X143Y128_DQ),
.I3(CLBLM_L_X92Y129_SLICE_X145Y129_A5Q),
.I4(CLBLM_L_X92Y129_SLICE_X145Y129_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y129_SLICE_X145Y129_DO5),
.O6(CLBLM_L_X92Y129_SLICE_X145Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y129_SLICE_X145Y129_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y129_SLICE_X145Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y129_SLICE_X145Y129_CO5),
.O6(CLBLM_L_X92Y129_SLICE_X145Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acccc0000)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_BLUT (
.I0(CLBLM_L_X92Y129_SLICE_X145Y129_AQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y129_SLICE_X145Y129_A5Q),
.I3(CLBLM_L_X92Y129_SLICE_X145Y129_CQ),
.I4(CLBLM_L_X92Y129_SLICE_X145Y129_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y129_SLICE_X145Y129_BO5),
.O6(CLBLM_L_X92Y129_SLICE_X145Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb800ff00b8000000)
  ) CLBLM_L_X92Y129_SLICE_X145Y129_ALUT (
.I0(CLBLM_R_X93Y129_SLICE_X146Y129_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X92Y129_SLICE_X145Y129_BO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X95Y131_SLICE_X150Y131_DO6),
.O5(CLBLM_L_X92Y129_SLICE_X145Y129_AO5),
.O6(CLBLM_L_X92Y129_SLICE_X145Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X144Y131_AO5),
.Q(CLBLM_L_X92Y131_SLICE_X144Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X144Y131_BO5),
.Q(CLBLM_L_X92Y131_SLICE_X144Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X144Y131_CO5),
.Q(CLBLM_L_X92Y131_SLICE_X144Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X144Y131_AO6),
.Q(CLBLM_L_X92Y131_SLICE_X144Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X144Y131_BO6),
.Q(CLBLM_L_X92Y131_SLICE_X144Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X144Y131_CO6),
.Q(CLBLM_L_X92Y131_SLICE_X144Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_DLUT (
.I0(CLBLM_L_X92Y131_SLICE_X145Y131_AQ),
.I1(CLBLM_L_X92Y131_SLICE_X145Y131_A5Q),
.I2(CLBLM_L_X92Y131_SLICE_X144Y131_AQ),
.I3(CLBLM_L_X92Y131_SLICE_X144Y131_A5Q),
.I4(CLBLM_L_X92Y131_SLICE_X144Y131_BQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y131_SLICE_X144Y131_DO5),
.O6(CLBLM_L_X92Y131_SLICE_X144Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00a0a88228822)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y131_SLICE_X144Y131_CQ),
.I2(CLBLM_R_X89Y130_SLICE_X140Y130_AQ),
.I3(CLBLM_R_X89Y128_SLICE_X140Y128_A5Q),
.I4(CLBLM_L_X92Y131_SLICE_X144Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y131_SLICE_X144Y131_CO5),
.O6(CLBLM_L_X92Y131_SLICE_X144Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00cc00c88884444)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_BLUT (
.I0(CLBLM_L_X90Y131_SLICE_X142Y131_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X90Y128_SLICE_X143Y128_D5Q),
.I3(CLBLM_L_X90Y130_SLICE_X142Y130_B5Q),
.I4(CLBLM_L_X92Y131_SLICE_X144Y131_BQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y131_SLICE_X144Y131_BO5),
.O6(CLBLM_L_X92Y131_SLICE_X144Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_L_X92Y131_SLICE_X144Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X92Y131_SLICE_X144Y131_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y131_SLICE_X145Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y131_SLICE_X144Y131_AO5),
.O6(CLBLM_L_X92Y131_SLICE_X144Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X145Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X145Y131_BO5),
.Q(CLBLM_L_X92Y131_SLICE_X145Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y131_SLICE_X145Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y131_SLICE_X145Y131_AO6),
.Q(CLBLM_L_X92Y131_SLICE_X145Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y131_SLICE_X145Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y131_SLICE_X145Y131_DO5),
.O6(CLBLM_L_X92Y131_SLICE_X145Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y131_SLICE_X145Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y131_SLICE_X145Y131_CO5),
.O6(CLBLM_L_X92Y131_SLICE_X145Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_L_X92Y131_SLICE_X145Y131_BLUT (
.I0(CLBLM_L_X92Y131_SLICE_X144Y131_A5Q),
.I1(CLBLM_L_X92Y131_SLICE_X145Y131_A5Q),
.I2(CLBLM_L_X92Y131_SLICE_X145Y131_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y131_SLICE_X144Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y131_SLICE_X145Y131_BO5),
.O6(CLBLM_L_X92Y131_SLICE_X145Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf300c000bb008800)
  ) CLBLM_L_X92Y131_SLICE_X145Y131_ALUT (
.I0(CLBLM_L_X92Y131_SLICE_X145Y131_BO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X93Y130_SLICE_X146Y130_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X97Y131_SLICE_X152Y131_CO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X92Y131_SLICE_X145Y131_AO5),
.O6(CLBLM_L_X92Y131_SLICE_X145Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y132_SLICE_X144Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y132_SLICE_X144Y132_DO5),
.O6(CLBLM_L_X92Y132_SLICE_X144Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y132_SLICE_X144Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y132_SLICE_X144Y132_CO5),
.O6(CLBLM_L_X92Y132_SLICE_X144Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y132_SLICE_X144Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y132_SLICE_X144Y132_BO5),
.O6(CLBLM_L_X92Y132_SLICE_X144Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X92Y132_SLICE_X144Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X92Y132_SLICE_X144Y132_AO5),
.O6(CLBLM_L_X92Y132_SLICE_X144Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y132_SLICE_X145Y132_BO5),
.Q(CLBLM_L_X92Y132_SLICE_X145Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y132_SLICE_X145Y132_CO5),
.Q(CLBLM_L_X92Y132_SLICE_X145Y132_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y132_SLICE_X145Y132_AO6),
.Q(CLBLM_L_X92Y132_SLICE_X145Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X92Y132_SLICE_X145Y132_CO6),
.Q(CLBLM_L_X92Y132_SLICE_X145Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_DLUT (
.I0(CLBLM_L_X92Y132_SLICE_X145Y132_C5Q),
.I1(CLBLM_L_X92Y132_SLICE_X145Y132_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y132_SLICE_X145Y132_A5Q),
.I4(CLBLM_L_X92Y132_SLICE_X145Y132_AQ),
.I5(CLBLM_L_X92Y131_SLICE_X144Y131_CQ),
.O5(CLBLM_L_X92Y132_SLICE_X145Y132_DO5),
.O6(CLBLM_L_X92Y132_SLICE_X145Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_CLUT (
.I0(CLBLM_L_X92Y132_SLICE_X145Y132_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y132_SLICE_X145Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X92Y132_SLICE_X145Y132_CO5),
.O6(CLBLM_L_X92Y132_SLICE_X145Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_BLUT (
.I0(CLBLM_L_X92Y132_SLICE_X145Y132_AQ),
.I1(CLBLM_L_X92Y132_SLICE_X145Y132_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y132_SLICE_X145Y132_CQ),
.I4(CLBLM_L_X92Y132_SLICE_X145Y132_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X92Y132_SLICE_X145Y132_BO5),
.O6(CLBLM_L_X92Y132_SLICE_X145Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ee2200000000)
  ) CLBLM_L_X92Y132_SLICE_X145Y132_ALUT (
.I0(CLBLM_R_X95Y132_SLICE_X150Y132_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X93Y132_SLICE_X146Y132_AQ),
.I3(CLBLM_L_X92Y132_SLICE_X145Y132_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X92Y132_SLICE_X145Y132_AO5),
.O6(CLBLM_L_X92Y132_SLICE_X145Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y111_SLICE_X148Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y111_SLICE_X148Y111_DO5),
.O6(CLBLM_L_X94Y111_SLICE_X148Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y111_SLICE_X148Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y111_SLICE_X148Y111_CO5),
.O6(CLBLM_L_X94Y111_SLICE_X148Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y111_SLICE_X148Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y111_SLICE_X148Y111_BO5),
.O6(CLBLM_L_X94Y111_SLICE_X148Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y111_SLICE_X148Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y111_SLICE_X148Y111_AO5),
.O6(CLBLM_L_X94Y111_SLICE_X148Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y111_SLICE_X149Y111_AO5),
.Q(CLBLM_L_X94Y111_SLICE_X149Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y111_SLICE_X149Y111_BO5),
.Q(CLBLM_L_X94Y111_SLICE_X149Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y111_SLICE_X149Y111_AO6),
.Q(CLBLM_L_X94Y111_SLICE_X149Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y111_SLICE_X149Y111_BO6),
.Q(CLBLM_L_X94Y111_SLICE_X149Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_DLUT (
.I0(CLBLM_L_X94Y111_SLICE_X149Y111_BQ),
.I1(CLBLM_R_X95Y111_SLICE_X150Y111_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X94Y111_SLICE_X149Y111_AQ),
.I4(CLBLM_L_X94Y111_SLICE_X149Y111_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X94Y111_SLICE_X149Y111_DO5),
.O6(CLBLM_L_X94Y111_SLICE_X149Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff550033f033f0)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_CLUT (
.I0(CLBLM_L_X94Y112_SLICE_X149Y112_A5Q),
.I1(CLBLM_R_X97Y111_SLICE_X152Y111_A5Q),
.I2(CLBLM_R_X93Y112_SLICE_X147Y112_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y111_SLICE_X149Y111_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X94Y111_SLICE_X149Y111_CO5),
.O6(CLBLM_L_X94Y111_SLICE_X149Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X94Y111_SLICE_X149Y111_AQ),
.I3(1'b1),
.I4(CLBLM_L_X94Y111_SLICE_X149Y111_BQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y111_SLICE_X149Y111_BO5),
.O6(CLBLM_L_X94Y111_SLICE_X149Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00a500a500)
  ) CLBLM_L_X94Y111_SLICE_X149Y111_ALUT (
.I0(CLBLM_R_X95Y113_SLICE_X150Y113_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X93Y114_SLICE_X147Y114_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y111_SLICE_X149Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y111_SLICE_X149Y111_AO5),
.O6(CLBLM_L_X94Y111_SLICE_X149Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X148Y112_AO5),
.Q(CLBLM_L_X94Y112_SLICE_X148Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X148Y112_BO5),
.Q(CLBLM_L_X94Y112_SLICE_X148Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X148Y112_AO6),
.Q(CLBLM_L_X94Y112_SLICE_X148Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X148Y112_BO6),
.Q(CLBLM_L_X94Y112_SLICE_X148Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55335533fff000f0)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_DLUT (
.I0(CLBLM_L_X94Y112_SLICE_X148Y112_A5Q),
.I1(CLBLM_R_X95Y112_SLICE_X150Y112_B5Q),
.I2(CLBLM_R_X93Y113_SLICE_X147Y113_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X93Y112_SLICE_X146Y112_CO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y112_SLICE_X148Y112_DO5),
.O6(CLBLM_L_X94Y112_SLICE_X148Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f3333ff00aaaa)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_CLUT (
.I0(CLBLM_R_X93Y112_SLICE_X146Y112_DO6),
.I1(CLBLM_R_X95Y112_SLICE_X150Y112_A5Q),
.I2(CLBLM_L_X94Y112_SLICE_X148Y112_AQ),
.I3(CLBLM_R_X93Y111_SLICE_X147Y111_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y112_SLICE_X148Y112_CO5),
.O6(CLBLM_L_X94Y112_SLICE_X148Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500c300c300)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_BLUT (
.I0(CLBLM_L_X94Y112_SLICE_X148Y112_DO6),
.I1(CLBLM_R_X93Y113_SLICE_X147Y113_A5Q),
.I2(CLBLM_L_X94Y112_SLICE_X149Y112_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y112_SLICE_X148Y112_BO5),
.O6(CLBLM_L_X94Y112_SLICE_X148Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_L_X94Y112_SLICE_X148Y112_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y112_SLICE_X148Y112_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y112_SLICE_X149Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y112_SLICE_X148Y112_AO5),
.O6(CLBLM_L_X94Y112_SLICE_X148Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X149Y112_AO5),
.Q(CLBLM_L_X94Y112_SLICE_X149Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X149Y112_BO5),
.Q(CLBLM_L_X94Y112_SLICE_X149Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X149Y112_AO6),
.Q(CLBLM_L_X94Y112_SLICE_X149Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y112_SLICE_X149Y112_BO6),
.Q(CLBLM_L_X94Y112_SLICE_X149Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y112_SLICE_X149Y112_DO5),
.O6(CLBLM_L_X94Y112_SLICE_X149Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32761054bafe98dc)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X94Y114_SLICE_X148Y114_CO6),
.I3(CLBLM_R_X95Y111_SLICE_X150Y111_A5Q),
.I4(CLBLM_R_X95Y111_SLICE_X150Y111_DO6),
.I5(CLBLM_L_X94Y112_SLICE_X149Y112_AQ),
.O5(CLBLM_L_X94Y112_SLICE_X149Y112_CO5),
.O6(CLBLM_L_X94Y112_SLICE_X149Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X94Y111_SLICE_X149Y111_A5Q),
.I4(CLBLM_L_X94Y112_SLICE_X149Y112_CO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y112_SLICE_X149Y112_BO5),
.O6(CLBLM_L_X94Y112_SLICE_X149Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cc00cc00)
  ) CLBLM_L_X94Y112_SLICE_X149Y112_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X95Y113_SLICE_X151Y113_AQ),
.I4(CLBLM_L_X94Y112_SLICE_X149Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y112_SLICE_X149Y112_AO5),
.O6(CLBLM_L_X94Y112_SLICE_X149Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y113_SLICE_X148Y113_AO5),
.Q(CLBLM_L_X94Y113_SLICE_X148Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y113_SLICE_X148Y113_BO5),
.Q(CLBLM_L_X94Y113_SLICE_X148Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y113_SLICE_X148Y113_AO6),
.Q(CLBLM_L_X94Y113_SLICE_X148Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y113_SLICE_X148Y113_BO6),
.Q(CLBLM_L_X94Y113_SLICE_X148Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c0f5cff5c005cf0)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_DLUT (
.I0(CLBLM_L_X94Y114_SLICE_X148Y114_AQ),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X94Y112_SLICE_X149Y112_B5Q),
.I5(CLBLM_L_X94Y117_SLICE_X148Y117_DO6),
.O5(CLBLM_L_X94Y113_SLICE_X148Y113_DO5),
.O6(CLBLM_L_X94Y113_SLICE_X148Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h454fe5ef404ae0ea)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X94Y114_SLICE_X148Y114_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y112_SLICE_X148Y112_B5Q),
.I4(CLBLM_L_X94Y113_SLICE_X148Y113_B5Q),
.I5(CLBLM_L_X94Y116_SLICE_X148Y116_DO6),
.O5(CLBLM_L_X94Y113_SLICE_X148Y113_CO5),
.O6(CLBLM_L_X94Y113_SLICE_X148Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888c0c0c0c0)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_BLUT (
.I0(CLBLM_L_X94Y113_SLICE_X148Y113_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X94Y114_SLICE_X148Y114_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y113_SLICE_X148Y113_BO5),
.O6(CLBLM_L_X94Y113_SLICE_X148Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500c300c300)
  ) CLBLM_L_X94Y113_SLICE_X148Y113_ALUT (
.I0(CLBLM_L_X94Y114_SLICE_X149Y114_CO6),
.I1(CLBLM_L_X92Y113_SLICE_X144Y113_A5Q),
.I2(CLBLM_R_X95Y112_SLICE_X150Y112_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y113_SLICE_X148Y113_AO5),
.O6(CLBLM_L_X94Y113_SLICE_X148Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y113_SLICE_X149Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y113_SLICE_X149Y113_AO5),
.Q(CLBLM_L_X94Y113_SLICE_X149Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y113_SLICE_X149Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y113_SLICE_X149Y113_AO6),
.Q(CLBLM_L_X94Y113_SLICE_X149Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y113_SLICE_X149Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y113_SLICE_X149Y113_DO5),
.O6(CLBLM_L_X94Y113_SLICE_X149Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_L_X94Y113_SLICE_X149Y113_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y114_SLICE_X150Y114_BQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y113_SLICE_X149Y113_A5Q),
.I4(CLBLM_L_X94Y113_SLICE_X149Y113_AQ),
.I5(CLBLM_L_X94Y114_SLICE_X149Y114_BQ),
.O5(CLBLM_L_X94Y113_SLICE_X149Y113_CO5),
.O6(CLBLM_L_X94Y113_SLICE_X149Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h47ff47cc47334700)
  ) CLBLM_L_X94Y113_SLICE_X149Y113_BLUT (
.I0(CLBLM_L_X94Y116_SLICE_X149Y116_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X95Y113_SLICE_X150Y113_B5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y115_SLICE_X149Y115_DO6),
.I5(CLBLM_L_X94Y113_SLICE_X149Y113_CO6),
.O5(CLBLM_L_X94Y113_SLICE_X149Y113_BO5),
.O6(CLBLM_L_X94Y113_SLICE_X149Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_L_X94Y113_SLICE_X149Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y114_SLICE_X150Y114_BQ),
.I2(CLBLM_L_X94Y113_SLICE_X149Y113_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y113_SLICE_X149Y113_AO5),
.O6(CLBLM_L_X94Y113_SLICE_X149Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X148Y114_AO5),
.Q(CLBLM_L_X94Y114_SLICE_X148Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X148Y114_BO5),
.Q(CLBLM_L_X94Y114_SLICE_X148Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X148Y114_AO6),
.Q(CLBLM_L_X94Y114_SLICE_X148Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X148Y114_BO6),
.Q(CLBLM_L_X94Y114_SLICE_X148Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y114_SLICE_X148Y114_DO5),
.O6(CLBLM_L_X94Y114_SLICE_X148Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_CLUT (
.I0(CLBLM_L_X94Y114_SLICE_X148Y114_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y113_SLICE_X147Y113_A5Q),
.I4(CLBLM_L_X94Y114_SLICE_X148Y114_B5Q),
.I5(CLBLM_L_X94Y115_SLICE_X148Y115_BQ),
.O5(CLBLM_L_X94Y114_SLICE_X148Y114_CO5),
.O6(CLBLM_L_X94Y114_SLICE_X148Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y114_SLICE_X148Y114_BQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y115_SLICE_X148Y115_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X94Y114_SLICE_X148Y114_BO5),
.O6(CLBLM_L_X94Y114_SLICE_X148Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ff000000)
  ) CLBLM_L_X94Y114_SLICE_X148Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y114_SLICE_X148Y114_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X94Y116_SLICE_X149Y116_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X94Y114_SLICE_X148Y114_AO5),
.O6(CLBLM_L_X94Y114_SLICE_X148Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X149Y114_AO5),
.Q(CLBLM_L_X94Y114_SLICE_X149Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X149Y114_BO5),
.Q(CLBLM_L_X94Y114_SLICE_X149Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X149Y114_AO6),
.Q(CLBLM_L_X94Y114_SLICE_X149Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y114_SLICE_X149Y114_BO6),
.Q(CLBLM_L_X94Y114_SLICE_X149Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33335555f0f0ff00)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_DLUT (
.I0(CLBLM_L_X94Y111_SLICE_X149Y111_A5Q),
.I1(CLBLM_L_X94Y114_SLICE_X148Y114_A5Q),
.I2(CLBLM_R_X93Y114_SLICE_X147Y114_CO6),
.I3(CLBLM_L_X94Y117_SLICE_X149Y117_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y114_SLICE_X149Y114_DO5),
.O6(CLBLM_L_X94Y114_SLICE_X149Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f00fffcacacaca)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_CLUT (
.I0(CLBLM_L_X92Y113_SLICE_X144Y113_CO6),
.I1(CLBLM_R_X95Y116_SLICE_X150Y116_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y114_SLICE_X149Y114_A5Q),
.I4(CLBLM_L_X98Y114_SLICE_X154Y114_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y114_SLICE_X149Y114_CO5),
.O6(CLBLM_L_X94Y114_SLICE_X149Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303000f000f0)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y113_SLICE_X149Y113_BO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X94Y115_SLICE_X149Y115_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y114_SLICE_X149Y114_BO5),
.O6(CLBLM_L_X94Y114_SLICE_X149Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X94Y114_SLICE_X149Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y114_SLICE_X149Y114_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y113_SLICE_X150Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y114_SLICE_X149Y114_AO5),
.O6(CLBLM_L_X94Y114_SLICE_X149Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X148Y115_AO5),
.Q(CLBLM_L_X94Y115_SLICE_X148Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X148Y115_BO5),
.Q(CLBLM_L_X94Y115_SLICE_X148Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X148Y115_CO5),
.Q(CLBLM_L_X94Y115_SLICE_X148Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X148Y115_AO6),
.Q(CLBLM_L_X94Y115_SLICE_X148Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X148Y115_BO6),
.Q(CLBLM_L_X94Y115_SLICE_X148Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X148Y115_CO6),
.Q(CLBLM_L_X94Y115_SLICE_X148Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_DLUT (
.I0(CLBLM_R_X95Y115_SLICE_X150Y115_AQ),
.I1(1'b1),
.I2(CLBLM_L_X94Y115_SLICE_X148Y115_AQ),
.I3(CLBLM_L_X94Y115_SLICE_X148Y115_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X93Y115_SLICE_X147Y115_AQ),
.O5(CLBLM_L_X94Y115_SLICE_X148Y115_DO5),
.O6(CLBLM_L_X94Y115_SLICE_X148Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00cc003300)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y115_SLICE_X149Y115_A5Q),
.I2(CLBLM_L_X94Y113_SLICE_X148Y113_DO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y117_SLICE_X149Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y115_SLICE_X148Y115_CO5),
.O6(CLBLM_L_X94Y115_SLICE_X148Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaa0a00a0a)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X94Y117_SLICE_X148Y117_A5Q),
.I3(CLBLM_L_X94Y113_SLICE_X148Y113_CO6),
.I4(CLBLM_L_X94Y115_SLICE_X148Y115_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y115_SLICE_X148Y115_BO5),
.O6(CLBLM_L_X94Y115_SLICE_X148Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_L_X94Y115_SLICE_X148Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X94Y115_SLICE_X148Y115_AQ),
.I3(CLBLM_R_X95Y115_SLICE_X150Y115_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y115_SLICE_X148Y115_AO5),
.O6(CLBLM_L_X94Y115_SLICE_X148Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X149Y115_AO5),
.Q(CLBLM_L_X94Y115_SLICE_X149Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X149Y115_BO5),
.Q(CLBLM_L_X94Y115_SLICE_X149Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X149Y115_AO6),
.Q(CLBLM_L_X94Y115_SLICE_X149Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y115_SLICE_X149Y115_BO6),
.Q(CLBLM_L_X94Y115_SLICE_X149Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_DLUT (
.I0(CLBLM_L_X94Y116_SLICE_X149Y116_C5Q),
.I1(CLBLM_L_X94Y114_SLICE_X149Y114_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X94Y115_SLICE_X149Y115_BQ),
.I4(CLBLM_L_X94Y115_SLICE_X149Y115_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X94Y115_SLICE_X149Y115_DO5),
.O6(CLBLM_L_X94Y115_SLICE_X149Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h757f252f707a202a)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X94Y117_SLICE_X149Y117_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y115_SLICE_X149Y115_A5Q),
.I4(CLBLM_L_X94Y115_SLICE_X149Y115_DO6),
.I5(CLBLM_R_X101Y121_SLICE_X159Y121_DO6),
.O5(CLBLM_L_X94Y115_SLICE_X149Y115_CO5),
.O6(CLBLM_L_X94Y115_SLICE_X149Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y115_SLICE_X149Y115_BQ),
.I2(CLBLM_L_X94Y114_SLICE_X149Y114_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y115_SLICE_X149Y115_BO5),
.O6(CLBLM_L_X94Y115_SLICE_X149Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_L_X94Y115_SLICE_X149Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y121_SLICE_X150Y121_A5Q),
.I2(CLBLM_L_X94Y116_SLICE_X149Y116_C5Q),
.I3(CLBLM_L_X94Y114_SLICE_X149Y114_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y115_SLICE_X149Y115_AO5),
.O6(CLBLM_L_X94Y115_SLICE_X149Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X148Y116_AO5),
.Q(CLBLM_L_X94Y116_SLICE_X148Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X148Y116_BO5),
.Q(CLBLM_L_X94Y116_SLICE_X148Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X148Y116_AO6),
.Q(CLBLM_L_X94Y116_SLICE_X148Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X148Y116_BO6),
.Q(CLBLM_L_X94Y116_SLICE_X148Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_DLUT (
.I0(CLBLM_R_X95Y118_SLICE_X150Y118_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y116_SLICE_X148Y116_BQ),
.I4(CLBLM_L_X94Y116_SLICE_X148Y116_B5Q),
.I5(CLBLM_L_X94Y117_SLICE_X148Y117_AQ),
.O5(CLBLM_L_X94Y116_SLICE_X148Y116_DO5),
.O6(CLBLM_L_X94Y116_SLICE_X148Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y116_SLICE_X148Y116_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y116_SLICE_X148Y116_A5Q),
.I4(CLBLM_R_X93Y116_SLICE_X147Y116_A5Q),
.I5(CLBLM_L_X94Y120_SLICE_X149Y120_BQ),
.O5(CLBLM_L_X94Y116_SLICE_X148Y116_CO5),
.O6(CLBLM_L_X94Y116_SLICE_X148Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y116_SLICE_X148Y116_BQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y117_SLICE_X148Y117_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y116_SLICE_X148Y116_BO5),
.O6(CLBLM_L_X94Y116_SLICE_X148Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_L_X94Y116_SLICE_X148Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X94Y116_SLICE_X148Y116_AQ),
.I3(CLBLM_L_X94Y120_SLICE_X149Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y116_SLICE_X148Y116_AO5),
.O6(CLBLM_L_X94Y116_SLICE_X148Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X149Y116_AO5),
.Q(CLBLM_L_X94Y116_SLICE_X149Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X149Y116_BO5),
.Q(CLBLM_L_X94Y116_SLICE_X149Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X149Y116_CO5),
.Q(CLBLM_L_X94Y116_SLICE_X149Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X149Y116_AO6),
.Q(CLBLM_L_X94Y116_SLICE_X149Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X149Y116_BO6),
.Q(CLBLM_L_X94Y116_SLICE_X149Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y116_SLICE_X149Y116_CO6),
.Q(CLBLM_L_X94Y116_SLICE_X149Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y116_SLICE_X149Y116_DO5),
.O6(CLBLM_L_X94Y116_SLICE_X149Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y115_SLICE_X149Y115_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y117_SLICE_X150Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y116_SLICE_X149Y116_CO5),
.O6(CLBLM_L_X94Y116_SLICE_X149Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y120_SLICE_X148Y120_AQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y116_SLICE_X149Y116_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y116_SLICE_X149Y116_BO5),
.O6(CLBLM_L_X94Y116_SLICE_X149Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLM_L_X94Y116_SLICE_X149Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y115_SLICE_X152Y115_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X93Y116_SLICE_X146Y116_A5Q),
.I4(CLBLM_L_X98Y117_SLICE_X155Y117_CO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y116_SLICE_X149Y116_AO5),
.O6(CLBLM_L_X94Y116_SLICE_X149Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X148Y117_AO5),
.Q(CLBLM_L_X94Y117_SLICE_X148Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X148Y117_BO5),
.Q(CLBLM_L_X94Y117_SLICE_X148Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X148Y117_AO6),
.Q(CLBLM_L_X94Y117_SLICE_X148Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X148Y117_BO6),
.Q(CLBLM_L_X94Y117_SLICE_X148Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_DLUT (
.I0(CLBLM_L_X94Y117_SLICE_X148Y117_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y117_SLICE_X148Y117_A5Q),
.I4(CLBLM_L_X94Y117_SLICE_X148Y117_B5Q),
.I5(CLBLM_R_X95Y118_SLICE_X150Y118_BQ),
.O5(CLBLM_L_X94Y117_SLICE_X148Y117_DO5),
.O6(CLBLM_L_X94Y117_SLICE_X148Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h777722225f0a5f0a)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X94Y118_SLICE_X148Y118_A5Q),
.I2(CLBLM_L_X94Y115_SLICE_X148Y115_B5Q),
.I3(CLBLM_R_X95Y118_SLICE_X151Y118_CO6),
.I4(CLBLM_L_X94Y117_SLICE_X148Y117_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X94Y117_SLICE_X148Y117_CO5),
.O6(CLBLM_L_X94Y117_SLICE_X148Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y117_SLICE_X148Y117_BQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y118_SLICE_X150Y118_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y117_SLICE_X148Y117_BO5),
.O6(CLBLM_L_X94Y117_SLICE_X148Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X94Y117_SLICE_X148Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y118_SLICE_X150Y118_AQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y117_SLICE_X148Y117_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y117_SLICE_X148Y117_AO5),
.O6(CLBLM_L_X94Y117_SLICE_X148Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X149Y117_AO5),
.Q(CLBLM_L_X94Y117_SLICE_X149Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X149Y117_BO5),
.Q(CLBLM_L_X94Y117_SLICE_X149Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X149Y117_AO6),
.Q(CLBLM_L_X94Y117_SLICE_X149Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y117_SLICE_X149Y117_BO6),
.Q(CLBLM_L_X94Y117_SLICE_X149Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_DLUT (
.I0(CLBLM_L_X94Y117_SLICE_X149Y117_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y117_SLICE_X150Y117_AQ),
.I4(CLBLM_L_X94Y117_SLICE_X149Y117_B5Q),
.I5(CLBLM_L_X94Y116_SLICE_X149Y116_CQ),
.O5(CLBLM_L_X94Y117_SLICE_X149Y117_DO5),
.O6(CLBLM_L_X94Y117_SLICE_X149Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h35353535fff00f00)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_CLUT (
.I0(CLBLM_L_X94Y115_SLICE_X148Y115_C5Q),
.I1(CLBLM_L_X94Y117_SLICE_X149Y117_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y117_SLICE_X150Y117_DO6),
.I4(CLBLM_L_X94Y117_SLICE_X149Y117_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y117_SLICE_X149Y117_CO5),
.O6(CLBLM_L_X94Y117_SLICE_X149Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y117_SLICE_X149Y117_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X94Y116_SLICE_X149Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y117_SLICE_X149Y117_BO5),
.O6(CLBLM_L_X94Y117_SLICE_X149Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X94Y117_SLICE_X149Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y117_SLICE_X149Y117_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X95Y120_SLICE_X150Y120_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y117_SLICE_X149Y117_AO5),
.O6(CLBLM_L_X94Y117_SLICE_X149Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y118_SLICE_X148Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y118_SLICE_X148Y118_AO5),
.Q(CLBLM_L_X94Y118_SLICE_X148Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y118_SLICE_X148Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y118_SLICE_X148Y118_AO6),
.Q(CLBLM_L_X94Y118_SLICE_X148Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y118_SLICE_X148Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y118_SLICE_X148Y118_DO5),
.O6(CLBLM_L_X94Y118_SLICE_X148Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y118_SLICE_X148Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y118_SLICE_X148Y118_CO5),
.O6(CLBLM_L_X94Y118_SLICE_X148Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00ccaa0fffccaa)
  ) CLBLM_L_X94Y118_SLICE_X148Y118_BLUT (
.I0(CLBLM_R_X97Y119_SLICE_X153Y119_DO6),
.I1(CLBLM_L_X94Y116_SLICE_X148Y116_DO6),
.I2(CLBLM_L_X94Y118_SLICE_X148Y118_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X93Y115_SLICE_X147Y115_B5Q),
.O5(CLBLM_L_X94Y118_SLICE_X148Y118_BO5),
.O6(CLBLM_L_X94Y118_SLICE_X148Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X94Y118_SLICE_X148Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y118_SLICE_X148Y118_A5Q),
.I2(CLBLM_L_X94Y117_SLICE_X149Y117_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y118_SLICE_X148Y118_AO5),
.O6(CLBLM_L_X94Y118_SLICE_X148Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y118_SLICE_X149Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y118_SLICE_X149Y118_AO5),
.Q(CLBLM_L_X94Y118_SLICE_X149Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y118_SLICE_X149Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y118_SLICE_X149Y118_AO6),
.Q(CLBLM_L_X94Y118_SLICE_X149Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y118_SLICE_X149Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y118_SLICE_X149Y118_DO5),
.O6(CLBLM_L_X94Y118_SLICE_X149Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y118_SLICE_X149Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y118_SLICE_X149Y118_CO5),
.O6(CLBLM_L_X94Y118_SLICE_X149Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e3e0232cefec2f2)
  ) CLBLM_L_X94Y118_SLICE_X149Y118_BLUT (
.I0(CLBLM_R_X95Y120_SLICE_X151Y120_CO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y114_SLICE_X146Y114_B5Q),
.I4(CLBLM_L_X94Y116_SLICE_X148Y116_CO6),
.I5(CLBLM_L_X94Y118_SLICE_X149Y118_A5Q),
.O5(CLBLM_L_X94Y118_SLICE_X149Y118_BO5),
.O6(CLBLM_L_X94Y118_SLICE_X149Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X94Y118_SLICE_X149Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y119_SLICE_X148Y119_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X94Y118_SLICE_X149Y118_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y118_SLICE_X149Y118_AO5),
.O6(CLBLM_L_X94Y118_SLICE_X149Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y119_SLICE_X148Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y119_SLICE_X148Y119_AO5),
.Q(CLBLM_L_X94Y119_SLICE_X148Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y119_SLICE_X148Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y119_SLICE_X148Y119_AO6),
.Q(CLBLM_L_X94Y119_SLICE_X148Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y119_SLICE_X148Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y119_SLICE_X148Y119_DO5),
.O6(CLBLM_L_X94Y119_SLICE_X148Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h330fffaa330f00aa)
  ) CLBLM_L_X94Y119_SLICE_X148Y119_CLUT (
.I0(CLBLM_R_X95Y121_SLICE_X151Y121_DO6),
.I1(CLBLM_L_X94Y119_SLICE_X148Y119_AQ),
.I2(CLBLM_R_X93Y115_SLICE_X146Y115_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X93Y118_SLICE_X147Y118_CO6),
.O5(CLBLM_L_X94Y119_SLICE_X148Y119_CO5),
.O6(CLBLM_L_X94Y119_SLICE_X148Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h23202f2ce3e0efec)
  ) CLBLM_L_X94Y119_SLICE_X148Y119_BLUT (
.I0(CLBLM_R_X93Y120_SLICE_X147Y120_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X97Y121_SLICE_X152Y121_DO6),
.I4(CLBLM_R_X93Y120_SLICE_X147Y120_C5Q),
.I5(CLBLM_L_X94Y120_SLICE_X148Y120_AQ),
.O5(CLBLM_L_X94Y119_SLICE_X148Y119_BO5),
.O6(CLBLM_L_X94Y119_SLICE_X148Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X94Y119_SLICE_X148Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y119_SLICE_X148Y119_A5Q),
.I2(CLBLM_L_X94Y118_SLICE_X148Y118_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y119_SLICE_X148Y119_AO5),
.O6(CLBLM_L_X94Y119_SLICE_X148Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y119_SLICE_X149Y119_AO5),
.Q(CLBLM_L_X94Y119_SLICE_X149Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y119_SLICE_X149Y119_BO5),
.Q(CLBLM_L_X94Y119_SLICE_X149Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y119_SLICE_X149Y119_AO6),
.Q(CLBLM_L_X94Y119_SLICE_X149Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y119_SLICE_X149Y119_BO6),
.Q(CLBLM_L_X94Y119_SLICE_X149Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_DLUT (
.I0(CLBLM_R_X95Y119_SLICE_X150Y119_AQ),
.I1(CLBLM_R_X93Y118_SLICE_X147Y118_A5Q),
.I2(CLBLM_L_X94Y119_SLICE_X149Y119_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X94Y119_SLICE_X149Y119_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y119_SLICE_X149Y119_DO5),
.O6(CLBLM_L_X94Y119_SLICE_X149Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0a300a3ffa30fa)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_CLUT (
.I0(CLBLM_R_X95Y119_SLICE_X150Y119_DO6),
.I1(CLBLM_L_X94Y119_SLICE_X148Y119_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X94Y119_SLICE_X149Y119_DO6),
.I5(CLBLM_R_X93Y115_SLICE_X146Y115_B5Q),
.O5(CLBLM_L_X94Y119_SLICE_X149Y119_CO5),
.O6(CLBLM_L_X94Y119_SLICE_X149Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_BLUT (
.I0(CLBLM_L_X94Y119_SLICE_X149Y119_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y119_SLICE_X150Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y119_SLICE_X149Y119_BO5),
.O6(CLBLM_L_X94Y119_SLICE_X149Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc84848484)
  ) CLBLM_L_X94Y119_SLICE_X149Y119_ALUT (
.I0(CLBLM_R_X95Y119_SLICE_X150Y119_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y119_SLICE_X150Y119_C5Q),
.I3(CLBLM_L_X94Y119_SLICE_X148Y119_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y119_SLICE_X149Y119_AO5),
.O6(CLBLM_L_X94Y119_SLICE_X149Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X148Y120_AO5),
.Q(CLBLM_L_X94Y120_SLICE_X148Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X148Y120_BO5),
.Q(CLBLM_L_X94Y120_SLICE_X148Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X148Y120_CO5),
.Q(CLBLM_L_X94Y120_SLICE_X148Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X148Y120_AO6),
.Q(CLBLM_L_X94Y120_SLICE_X148Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X148Y120_BO6),
.Q(CLBLM_L_X94Y120_SLICE_X148Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X148Y120_CO6),
.Q(CLBLM_L_X94Y120_SLICE_X148Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bbf5f511bba0a0)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y120_SLICE_X147Y120_CQ),
.I2(CLBLM_R_X93Y120_SLICE_X146Y120_DO6),
.I3(CLBLM_L_X94Y120_SLICE_X148Y120_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y120_SLICE_X150Y120_CO6),
.O5(CLBLM_L_X94Y120_SLICE_X148Y120_DO5),
.O6(CLBLM_L_X94Y120_SLICE_X148Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00c300c300)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y122_SLICE_X150Y122_B5Q),
.I2(CLBLM_R_X93Y124_SLICE_X147Y124_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y120_SLICE_X148Y120_DO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y120_SLICE_X148Y120_CO5),
.O6(CLBLM_L_X94Y120_SLICE_X148Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc88884444)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_BLUT (
.I0(CLBLM_R_X95Y120_SLICE_X150Y120_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_L_X94Y119_SLICE_X148Y119_BO6),
.I4(CLBLM_L_X94Y120_SLICE_X148Y120_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y120_SLICE_X148Y120_BO5),
.O6(CLBLM_L_X94Y120_SLICE_X148Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_L_X94Y120_SLICE_X148Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y120_SLICE_X148Y120_A5Q),
.I2(CLBLM_L_X92Y120_SLICE_X144Y120_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y120_SLICE_X148Y120_AO5),
.O6(CLBLM_L_X94Y120_SLICE_X148Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X149Y120_AO5),
.Q(CLBLM_L_X94Y120_SLICE_X149Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X149Y120_BO5),
.Q(CLBLM_L_X94Y120_SLICE_X149Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X149Y120_AO6),
.Q(CLBLM_L_X94Y120_SLICE_X149Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y120_SLICE_X149Y120_BO6),
.Q(CLBLM_L_X94Y120_SLICE_X149Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y120_SLICE_X149Y120_DO5),
.O6(CLBLM_L_X94Y120_SLICE_X149Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0add885f5fdd88)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y116_SLICE_X147Y116_CO6),
.I2(CLBLM_L_X94Y118_SLICE_X149Y118_AQ),
.I3(CLBLM_R_X95Y123_SLICE_X150Y123_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X93Y114_SLICE_X146Y114_A5Q),
.O5(CLBLM_L_X94Y120_SLICE_X149Y120_CO5),
.O6(CLBLM_L_X94Y120_SLICE_X149Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300aa005500)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_BLUT (
.I0(CLBLM_R_X95Y120_SLICE_X151Y120_A5Q),
.I1(CLBLM_L_X94Y118_SLICE_X149Y118_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y119_SLICE_X149Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y120_SLICE_X149Y120_BO5),
.O6(CLBLM_L_X94Y120_SLICE_X149Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00a500a500)
  ) CLBLM_L_X94Y120_SLICE_X149Y120_ALUT (
.I0(CLBLM_L_X94Y120_SLICE_X149Y120_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X95Y120_SLICE_X151Y120_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y120_SLICE_X149Y120_CO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y120_SLICE_X149Y120_AO5),
.O6(CLBLM_L_X94Y120_SLICE_X149Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y121_SLICE_X148Y121_BO5),
.Q(CLBLM_L_X94Y121_SLICE_X148Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y121_SLICE_X148Y121_CO5),
.Q(CLBLM_L_X94Y121_SLICE_X148Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y121_SLICE_X148Y121_AO6),
.Q(CLBLM_L_X94Y121_SLICE_X148Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y121_SLICE_X148Y121_CO6),
.Q(CLBLM_L_X94Y121_SLICE_X148Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X94Y121_SLICE_X148Y121_AQ),
.I2(CLBLM_R_X97Y120_SLICE_X153Y120_DQ),
.I3(CLBLM_L_X94Y121_SLICE_X148Y121_A5Q),
.I4(CLBLM_L_X94Y121_SLICE_X148Y121_CQ),
.I5(CLBLM_R_X93Y121_SLICE_X147Y121_C5Q),
.O5(CLBLM_L_X94Y121_SLICE_X148Y121_DO5),
.O6(CLBLM_L_X94Y121_SLICE_X148Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y121_SLICE_X148Y121_AQ),
.I2(1'b1),
.I3(CLBLM_L_X92Y120_SLICE_X145Y120_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y121_SLICE_X148Y121_CO5),
.O6(CLBLM_L_X94Y121_SLICE_X148Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996ff000000)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_BLUT (
.I0(CLBLM_L_X94Y121_SLICE_X148Y121_CQ),
.I1(CLBLM_L_X94Y121_SLICE_X148Y121_A5Q),
.I2(CLBLM_L_X94Y121_SLICE_X148Y121_AQ),
.I3(CLBLM_R_X93Y121_SLICE_X147Y121_C5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X94Y121_SLICE_X148Y121_BO5),
.O6(CLBLM_L_X94Y121_SLICE_X148Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heee200002e220000)
  ) CLBLM_L_X94Y121_SLICE_X148Y121_ALUT (
.I0(CLBLM_L_X90Y121_SLICE_X143Y121_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X94Y121_SLICE_X148Y121_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_L_X92Y119_SLICE_X145Y119_AQ),
.O5(CLBLM_L_X94Y121_SLICE_X148Y121_AO5),
.O6(CLBLM_L_X94Y121_SLICE_X148Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y121_SLICE_X149Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y121_SLICE_X149Y121_AO5),
.Q(CLBLM_L_X94Y121_SLICE_X149Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y121_SLICE_X149Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y121_SLICE_X149Y121_AO6),
.Q(CLBLM_L_X94Y121_SLICE_X149Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y121_SLICE_X149Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y121_SLICE_X149Y121_DO5),
.O6(CLBLM_L_X94Y121_SLICE_X149Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff33f0550033f0)
  ) CLBLM_L_X94Y121_SLICE_X149Y121_CLUT (
.I0(CLBLM_L_X94Y121_SLICE_X149Y121_A5Q),
.I1(CLBLM_R_X93Y119_SLICE_X146Y119_B5Q),
.I2(CLBLM_R_X95Y123_SLICE_X151Y123_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X93Y119_SLICE_X147Y119_CO6),
.O5(CLBLM_L_X94Y121_SLICE_X149Y121_CO5),
.O6(CLBLM_L_X94Y121_SLICE_X149Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d7f193b4c6e082a)
  ) CLBLM_L_X94Y121_SLICE_X149Y121_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X94Y121_SLICE_X149Y121_AQ),
.I3(CLBLM_R_X93Y119_SLICE_X146Y119_A5Q),
.I4(CLBLM_R_X93Y119_SLICE_X146Y119_DO6),
.I5(CLBLM_R_X95Y126_SLICE_X150Y126_CO6),
.O5(CLBLM_L_X94Y121_SLICE_X149Y121_BO5),
.O6(CLBLM_L_X94Y121_SLICE_X149Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000a0a0a0a0)
  ) CLBLM_L_X94Y121_SLICE_X149Y121_ALUT (
.I0(CLBLM_L_X94Y118_SLICE_X149Y118_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X94Y121_SLICE_X149Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y121_SLICE_X149Y121_AO5),
.O6(CLBLM_L_X94Y121_SLICE_X149Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_DO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_CO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_BO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X148Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X148Y122_AO5),
.O6(CLBLM_L_X94Y122_SLICE_X148Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y122_SLICE_X149Y122_AO5),
.Q(CLBLM_L_X94Y122_SLICE_X149Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y122_SLICE_X149Y122_BO5),
.Q(CLBLM_L_X94Y122_SLICE_X149Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y122_SLICE_X149Y122_AO6),
.Q(CLBLM_L_X94Y122_SLICE_X149Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y122_SLICE_X149Y122_BO6),
.Q(CLBLM_L_X94Y122_SLICE_X149Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_DO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_CO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00a500a500)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_BLUT (
.I0(CLBLM_R_X95Y123_SLICE_X150Y123_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X94Y120_SLICE_X149Y120_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y121_SLICE_X149Y121_CO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_BO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300aa005500)
  ) CLBLM_L_X94Y122_SLICE_X149Y122_ALUT (
.I0(CLBLM_L_X94Y122_SLICE_X149Y122_B5Q),
.I1(CLBLM_L_X94Y121_SLICE_X149Y121_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y123_SLICE_X151Y123_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y122_SLICE_X149Y122_AO5),
.O6(CLBLM_L_X94Y122_SLICE_X149Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y123_SLICE_X148Y123_BO5),
.Q(CLBLM_L_X94Y123_SLICE_X148Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y123_SLICE_X148Y123_CO5),
.Q(CLBLM_L_X94Y123_SLICE_X148Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y123_SLICE_X148Y123_AO6),
.Q(CLBLM_L_X94Y123_SLICE_X148Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y123_SLICE_X148Y123_CO6),
.Q(CLBLM_L_X94Y123_SLICE_X148Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_DLUT (
.I0(CLBLM_L_X94Y123_SLICE_X148Y123_C5Q),
.I1(CLBLM_L_X94Y123_SLICE_X148Y123_AQ),
.I2(CLBLM_L_X92Y122_SLICE_X144Y122_C5Q),
.I3(CLBLM_L_X94Y123_SLICE_X148Y123_A5Q),
.I4(CLBLM_L_X94Y123_SLICE_X148Y123_CQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y123_SLICE_X148Y123_DO5),
.O6(CLBLM_L_X94Y123_SLICE_X148Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X94Y123_SLICE_X148Y123_AQ),
.I3(1'b1),
.I4(CLBLM_L_X94Y123_SLICE_X148Y123_CQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y123_SLICE_X148Y123_CO5),
.O6(CLBLM_L_X94Y123_SLICE_X148Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_BLUT (
.I0(CLBLM_L_X94Y123_SLICE_X148Y123_CQ),
.I1(CLBLM_L_X94Y123_SLICE_X148Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X94Y123_SLICE_X148Y123_AQ),
.I4(CLBLM_L_X94Y123_SLICE_X148Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y123_SLICE_X148Y123_BO5),
.O6(CLBLM_L_X94Y123_SLICE_X148Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b0c08070304000)
  ) CLBLM_L_X94Y123_SLICE_X148Y123_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X94Y123_SLICE_X148Y123_BO6),
.I4(CLBLM_R_X95Y124_SLICE_X151Y124_DO6),
.I5(CLBLM_L_X94Y124_SLICE_X148Y124_A5Q),
.O5(CLBLM_L_X94Y123_SLICE_X148Y123_AO5),
.O6(CLBLM_L_X94Y123_SLICE_X148Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y123_SLICE_X149Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y123_SLICE_X149Y123_DO5),
.O6(CLBLM_L_X94Y123_SLICE_X149Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y123_SLICE_X149Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y123_SLICE_X149Y123_CO5),
.O6(CLBLM_L_X94Y123_SLICE_X149Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y123_SLICE_X149Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y123_SLICE_X149Y123_BO5),
.O6(CLBLM_L_X94Y123_SLICE_X149Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y123_SLICE_X149Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y123_SLICE_X149Y123_AO5),
.O6(CLBLM_L_X94Y123_SLICE_X149Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X148Y124_AO5),
.Q(CLBLM_L_X94Y124_SLICE_X148Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X148Y124_BO5),
.Q(CLBLM_L_X94Y124_SLICE_X148Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X148Y124_CO5),
.Q(CLBLM_L_X94Y124_SLICE_X148Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X148Y124_AO6),
.Q(CLBLM_L_X94Y124_SLICE_X148Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X148Y124_BO6),
.Q(CLBLM_L_X94Y124_SLICE_X148Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X148Y124_CO6),
.Q(CLBLM_L_X94Y124_SLICE_X148Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X94Y125_SLICE_X148Y125_BQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y124_SLICE_X148Y124_BQ),
.I4(CLBLM_L_X94Y124_SLICE_X148Y124_B5Q),
.I5(CLBLM_R_X93Y124_SLICE_X147Y124_B5Q),
.O5(CLBLM_L_X94Y124_SLICE_X148Y124_DO5),
.O6(CLBLM_L_X94Y124_SLICE_X148Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_CLUT (
.I0(CLBLM_L_X94Y123_SLICE_X148Y123_A5Q),
.I1(CLBLM_L_X94Y124_SLICE_X148Y124_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y125_SLICE_X147Y125_A5Q),
.I4(CLBLM_R_X93Y124_SLICE_X146Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y124_SLICE_X148Y124_CO5),
.O6(CLBLM_L_X94Y124_SLICE_X148Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_BLUT (
.I0(CLBLM_L_X94Y125_SLICE_X148Y125_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X94Y124_SLICE_X148Y124_BQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y124_SLICE_X148Y124_BO5),
.O6(CLBLM_L_X94Y124_SLICE_X148Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_L_X94Y124_SLICE_X148Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y124_SLICE_X148Y124_A5Q),
.I2(CLBLM_R_X93Y126_SLICE_X146Y126_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y124_SLICE_X148Y124_AO5),
.O6(CLBLM_L_X94Y124_SLICE_X148Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X149Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X149Y124_AO5),
.Q(CLBLM_L_X94Y124_SLICE_X149Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y124_SLICE_X149Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y124_SLICE_X149Y124_AO6),
.Q(CLBLM_L_X94Y124_SLICE_X149Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y124_SLICE_X149Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y124_SLICE_X149Y124_DO5),
.O6(CLBLM_L_X94Y124_SLICE_X149Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X94Y124_SLICE_X149Y124_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X94Y128_SLICE_X149Y128_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X94Y124_SLICE_X149Y124_A5Q),
.I4(CLBLM_L_X94Y124_SLICE_X149Y124_AQ),
.I5(CLBLM_L_X98Y128_SLICE_X154Y128_AQ),
.O5(CLBLM_L_X94Y124_SLICE_X149Y124_CO5),
.O6(CLBLM_L_X94Y124_SLICE_X149Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3077fc773044fc44)
  ) CLBLM_L_X94Y124_SLICE_X149Y124_BLUT (
.I0(CLBLM_R_X93Y124_SLICE_X147Y124_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X93Y124_SLICE_X147Y124_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X94Y124_SLICE_X148Y124_AQ),
.I5(CLBLM_L_X94Y124_SLICE_X149Y124_CO6),
.O5(CLBLM_L_X94Y124_SLICE_X149Y124_BO5),
.O6(CLBLM_L_X94Y124_SLICE_X149Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_L_X94Y124_SLICE_X149Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X94Y124_SLICE_X149Y124_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y128_SLICE_X154Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y124_SLICE_X149Y124_AO5),
.O6(CLBLM_L_X94Y124_SLICE_X149Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X148Y125_AO5),
.Q(CLBLM_L_X94Y125_SLICE_X148Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X148Y125_BO5),
.Q(CLBLM_L_X94Y125_SLICE_X148Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X148Y125_AO6),
.Q(CLBLM_L_X94Y125_SLICE_X148Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X148Y125_BO6),
.Q(CLBLM_L_X94Y125_SLICE_X148Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_DLUT (
.I0(CLBLM_L_X94Y125_SLICE_X149Y125_A5Q),
.I1(CLBLM_L_X94Y125_SLICE_X149Y125_AQ),
.I2(CLBLM_R_X93Y125_SLICE_X147Y125_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y125_SLICE_X149Y125_DQ),
.I5(CLBLM_L_X94Y125_SLICE_X149Y125_C5Q),
.O5(CLBLM_L_X94Y125_SLICE_X148Y125_DO5),
.O6(CLBLM_L_X94Y125_SLICE_X148Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff330055f055f0)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_CLUT (
.I0(CLBLM_R_X93Y120_SLICE_X146Y120_A5Q),
.I1(CLBLM_L_X94Y125_SLICE_X148Y125_AQ),
.I2(CLBLM_R_X95Y125_SLICE_X151Y125_CO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y124_SLICE_X148Y124_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X94Y125_SLICE_X148Y125_CO5),
.O6(CLBLM_L_X94Y125_SLICE_X148Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ccccc00cc00c)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X94Y122_SLICE_X149Y122_A5Q),
.I3(CLBLM_R_X95Y126_SLICE_X150Y126_A5Q),
.I4(CLBLM_L_X94Y125_SLICE_X148Y125_CO6),
.I5(1'b1),
.O5(CLBLM_L_X94Y125_SLICE_X148Y125_BO5),
.O6(CLBLM_L_X94Y125_SLICE_X148Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000000f000f00)
  ) CLBLM_L_X94Y125_SLICE_X148Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X94Y125_SLICE_X148Y125_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y121_SLICE_X149Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y125_SLICE_X148Y125_AO5),
.O6(CLBLM_L_X94Y125_SLICE_X148Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X149Y125_BO5),
.Q(CLBLM_L_X94Y125_SLICE_X149Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X149Y125_CO5),
.Q(CLBLM_L_X94Y125_SLICE_X149Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X149Y125_DO5),
.Q(CLBLM_L_X94Y125_SLICE_X149Y125_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X149Y125_AO6),
.Q(CLBLM_L_X94Y125_SLICE_X149Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X149Y125_CO6),
.Q(CLBLM_L_X94Y125_SLICE_X149Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y125_SLICE_X149Y125_DO6),
.Q(CLBLM_L_X94Y125_SLICE_X149Y125_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y128_SLICE_X150Y128_BQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y125_SLICE_X149Y125_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y125_SLICE_X149Y125_DO5),
.O6(CLBLM_L_X94Y125_SLICE_X149Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X94Y125_SLICE_X149Y125_DQ),
.I3(CLBLM_R_X95Y125_SLICE_X150Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y125_SLICE_X149Y125_CO5),
.O6(CLBLM_L_X94Y125_SLICE_X149Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acccc0000)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_BLUT (
.I0(CLBLM_L_X94Y125_SLICE_X149Y125_AQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X94Y125_SLICE_X149Y125_A5Q),
.I3(CLBLM_L_X94Y125_SLICE_X149Y125_DQ),
.I4(CLBLM_L_X94Y125_SLICE_X149Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y125_SLICE_X149Y125_BO5),
.O6(CLBLM_L_X94Y125_SLICE_X149Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee002200e200e200)
  ) CLBLM_L_X94Y125_SLICE_X149Y125_ALUT (
.I0(CLBLM_L_X98Y126_SLICE_X155Y126_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X94Y125_SLICE_X149Y125_BO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y127_SLICE_X149Y127_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X94Y125_SLICE_X149Y125_AO5),
.O6(CLBLM_L_X94Y125_SLICE_X149Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X148Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X148Y126_DO5),
.O6(CLBLM_L_X94Y126_SLICE_X148Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X148Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X148Y126_CO5),
.O6(CLBLM_L_X94Y126_SLICE_X148Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X148Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X148Y126_BO5),
.O6(CLBLM_L_X94Y126_SLICE_X148Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X148Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X148Y126_AO5),
.O6(CLBLM_L_X94Y126_SLICE_X148Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X149Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X149Y126_DO5),
.O6(CLBLM_L_X94Y126_SLICE_X149Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X149Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X149Y126_CO5),
.O6(CLBLM_L_X94Y126_SLICE_X149Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y126_SLICE_X149Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y126_SLICE_X149Y126_BO5),
.O6(CLBLM_L_X94Y126_SLICE_X149Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_L_X94Y126_SLICE_X149Y126_ALUT (
.I0(CLBLM_L_X94Y127_SLICE_X149Y127_B5Q),
.I1(CLBLM_L_X94Y125_SLICE_X149Y125_D5Q),
.I2(CLBLM_R_X93Y125_SLICE_X147Y125_AQ),
.I3(CLBLM_L_X94Y127_SLICE_X149Y127_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y128_SLICE_X150Y128_BQ),
.O5(CLBLM_L_X94Y126_SLICE_X149Y126_AO5),
.O6(CLBLM_L_X94Y126_SLICE_X149Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y127_SLICE_X148Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X148Y127_DO5),
.O6(CLBLM_L_X94Y127_SLICE_X148Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y127_SLICE_X148Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X148Y127_CO5),
.O6(CLBLM_L_X94Y127_SLICE_X148Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y127_SLICE_X148Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X148Y127_BO5),
.O6(CLBLM_L_X94Y127_SLICE_X148Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y127_SLICE_X148Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X148Y127_AO5),
.O6(CLBLM_L_X94Y127_SLICE_X148Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y127_SLICE_X149Y127_AO5),
.Q(CLBLM_L_X94Y127_SLICE_X149Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y127_SLICE_X149Y127_CO5),
.Q(CLBLM_L_X94Y127_SLICE_X149Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y127_SLICE_X149Y127_AO6),
.Q(CLBLM_L_X94Y127_SLICE_X149Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y127_SLICE_X149Y127_BO6),
.Q(CLBLM_L_X94Y127_SLICE_X149Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X149Y127_DO5),
.O6(CLBLM_L_X94Y127_SLICE_X149Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_CLUT (
.I0(CLBLM_L_X94Y125_SLICE_X149Y125_D5Q),
.I1(CLBLM_R_X95Y128_SLICE_X150Y128_BQ),
.I2(CLBLM_L_X94Y127_SLICE_X149Y127_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y127_SLICE_X149Y127_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X149Y127_CO5),
.O6(CLBLM_L_X94Y127_SLICE_X149Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heee222e200000000)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_BLUT (
.I0(CLBLM_R_X97Y126_SLICE_X153Y126_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X94Y127_SLICE_X149Y127_CO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y127_SLICE_X149Y127_A5Q),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X94Y127_SLICE_X149Y127_BO5),
.O6(CLBLM_L_X94Y127_SLICE_X149Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X94Y127_SLICE_X149Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y127_SLICE_X149Y127_A5Q),
.I2(CLBLM_L_X94Y130_SLICE_X149Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y127_SLICE_X149Y127_AO5),
.O6(CLBLM_L_X94Y127_SLICE_X149Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y128_SLICE_X148Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y128_SLICE_X148Y128_DO5),
.O6(CLBLM_L_X94Y128_SLICE_X148Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y128_SLICE_X148Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y128_SLICE_X148Y128_CO5),
.O6(CLBLM_L_X94Y128_SLICE_X148Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y128_SLICE_X148Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y128_SLICE_X148Y128_BO5),
.O6(CLBLM_L_X94Y128_SLICE_X148Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y128_SLICE_X148Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y128_SLICE_X148Y128_AO5),
.O6(CLBLM_L_X94Y128_SLICE_X148Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y128_SLICE_X149Y128_BO5),
.Q(CLBLM_L_X94Y128_SLICE_X149Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y128_SLICE_X149Y128_CO5),
.Q(CLBLM_L_X94Y128_SLICE_X149Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y128_SLICE_X149Y128_AO6),
.Q(CLBLM_L_X94Y128_SLICE_X149Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y128_SLICE_X149Y128_CO6),
.Q(CLBLM_L_X94Y128_SLICE_X149Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd8d88dd88d8dd8)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X93Y128_SLICE_X147Y128_DQ),
.I2(CLBLM_L_X94Y129_SLICE_X148Y129_B5Q),
.I3(CLBLM_L_X94Y128_SLICE_X149Y128_A5Q),
.I4(CLBLM_L_X94Y128_SLICE_X149Y128_AQ),
.I5(CLBLM_L_X94Y128_SLICE_X149Y128_CQ),
.O5(CLBLM_L_X94Y128_SLICE_X149Y128_DO5),
.O6(CLBLM_L_X94Y128_SLICE_X149Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cc00cc00)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_L_X94Y124_SLICE_X149Y124_A5Q),
.I4(CLBLM_L_X94Y128_SLICE_X149Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y128_SLICE_X149Y128_CO5),
.O6(CLBLM_L_X94Y128_SLICE_X149Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y128_SLICE_X149Y128_A5Q),
.I2(CLBLM_L_X94Y128_SLICE_X149Y128_AQ),
.I3(CLBLM_L_X94Y128_SLICE_X149Y128_CQ),
.I4(CLBLM_L_X94Y129_SLICE_X148Y129_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y128_SLICE_X149Y128_BO5),
.O6(CLBLM_L_X94Y128_SLICE_X149Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heee22e2200000000)
  ) CLBLM_L_X94Y128_SLICE_X149Y128_ALUT (
.I0(CLBLM_R_X97Y128_SLICE_X153Y128_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X94Y128_SLICE_X149Y128_BO6),
.I4(CLBLM_L_X94Y130_SLICE_X149Y130_AQ),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X94Y128_SLICE_X149Y128_AO5),
.O6(CLBLM_L_X94Y128_SLICE_X149Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y129_SLICE_X148Y129_BO5),
.Q(CLBLM_L_X94Y129_SLICE_X148Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y129_SLICE_X148Y129_AO5),
.Q(CLBLM_L_X94Y129_SLICE_X148Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y129_SLICE_X148Y129_BO6),
.Q(CLBLM_L_X94Y129_SLICE_X148Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X148Y129_DO5),
.O6(CLBLM_L_X94Y129_SLICE_X148Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_CLUT (
.I0(CLBLM_L_X94Y130_SLICE_X148Y130_AQ),
.I1(CLBLM_L_X94Y129_SLICE_X148Y129_AQ),
.I2(CLBLM_R_X95Y129_SLICE_X150Y129_C5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y129_SLICE_X148Y129_BQ),
.I5(CLBLM_R_X93Y128_SLICE_X147Y128_A5Q),
.O5(CLBLM_L_X94Y129_SLICE_X148Y129_CO5),
.O6(CLBLM_L_X94Y129_SLICE_X148Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y128_SLICE_X149Y128_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X94Y130_SLICE_X148Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X148Y129_BO5),
.O6(CLBLM_L_X94Y129_SLICE_X148Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f000f000)
  ) CLBLM_L_X94Y129_SLICE_X148Y129_ALUT (
.I0(CLBLM_L_X94Y129_SLICE_X148Y129_AQ),
.I1(CLBLM_L_X94Y129_SLICE_X148Y129_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y129_SLICE_X150Y129_C5Q),
.I4(CLBLM_L_X94Y130_SLICE_X148Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X148Y129_AO5),
.O6(CLBLM_L_X94Y129_SLICE_X148Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y129_SLICE_X149Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X149Y129_DO5),
.O6(CLBLM_L_X94Y129_SLICE_X149Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y129_SLICE_X149Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X149Y129_CO5),
.O6(CLBLM_L_X94Y129_SLICE_X149Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y129_SLICE_X149Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X149Y129_BO5),
.O6(CLBLM_L_X94Y129_SLICE_X149Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y129_SLICE_X149Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y129_SLICE_X149Y129_AO5),
.O6(CLBLM_L_X94Y129_SLICE_X149Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y130_SLICE_X148Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y130_SLICE_X148Y130_AO6),
.Q(CLBLM_L_X94Y130_SLICE_X148Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y130_SLICE_X148Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X148Y130_DO5),
.O6(CLBLM_L_X94Y130_SLICE_X148Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y130_SLICE_X148Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X148Y130_CO5),
.O6(CLBLM_L_X94Y130_SLICE_X148Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y130_SLICE_X148Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X148Y130_BO5),
.O6(CLBLM_L_X94Y130_SLICE_X148Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f0c0f0a000c000)
  ) CLBLM_L_X94Y130_SLICE_X148Y130_ALUT (
.I0(CLBLM_R_X95Y131_SLICE_X150Y131_A5Q),
.I1(CLBLM_L_X94Y129_SLICE_X148Y129_AO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X97Y130_SLICE_X152Y130_CO6),
.O5(CLBLM_L_X94Y130_SLICE_X148Y130_AO5),
.O6(CLBLM_L_X94Y130_SLICE_X148Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y130_SLICE_X149Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y130_SLICE_X149Y130_AO5),
.Q(CLBLM_L_X94Y130_SLICE_X149Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X94Y130_SLICE_X149Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X94Y130_SLICE_X149Y130_AO6),
.Q(CLBLM_L_X94Y130_SLICE_X149Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y130_SLICE_X149Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X149Y130_DO5),
.O6(CLBLM_L_X94Y130_SLICE_X149Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y130_SLICE_X149Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X149Y130_CO5),
.O6(CLBLM_L_X94Y130_SLICE_X149Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y130_SLICE_X149Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X149Y130_BO5),
.O6(CLBLM_L_X94Y130_SLICE_X149Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X94Y130_SLICE_X149Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y132_SLICE_X151Y132_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X94Y130_SLICE_X149Y130_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X94Y130_SLICE_X149Y130_AO5),
.O6(CLBLM_L_X94Y130_SLICE_X149Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X148Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X148Y132_DO5),
.O6(CLBLM_L_X94Y132_SLICE_X148Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X148Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X148Y132_CO5),
.O6(CLBLM_L_X94Y132_SLICE_X148Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X148Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X148Y132_BO5),
.O6(CLBLM_L_X94Y132_SLICE_X148Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X148Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X148Y132_AO5),
.O6(CLBLM_L_X94Y132_SLICE_X148Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X149Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X149Y132_DO5),
.O6(CLBLM_L_X94Y132_SLICE_X149Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X149Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X149Y132_CO5),
.O6(CLBLM_L_X94Y132_SLICE_X149Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X94Y132_SLICE_X149Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X94Y132_SLICE_X149Y132_BO5),
.O6(CLBLM_L_X94Y132_SLICE_X149Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69ff9600690096)
  ) CLBLM_L_X94Y132_SLICE_X149Y132_ALUT (
.I0(CLBLM_R_X95Y132_SLICE_X151Y132_CQ),
.I1(CLBLM_R_X95Y132_SLICE_X150Y132_C5Q),
.I2(CLBLM_R_X97Y132_SLICE_X152Y132_DQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X95Y132_SLICE_X151Y132_B5Q),
.I5(CLBLM_R_X93Y131_SLICE_X147Y131_A5Q),
.O5(CLBLM_L_X94Y132_SLICE_X149Y132_AO5),
.O6(CLBLM_L_X94Y132_SLICE_X149Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y110_SLICE_X154Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y110_SLICE_X154Y110_AO5),
.Q(CLBLM_L_X98Y110_SLICE_X154Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y110_SLICE_X154Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y110_SLICE_X154Y110_AO6),
.Q(CLBLM_L_X98Y110_SLICE_X154Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y110_SLICE_X154Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X154Y110_DO5),
.O6(CLBLM_L_X98Y110_SLICE_X154Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y110_SLICE_X154Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X154Y110_CO5),
.O6(CLBLM_L_X98Y110_SLICE_X154Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_L_X98Y110_SLICE_X154Y110_BLUT (
.I0(CLBLM_L_X98Y111_SLICE_X154Y111_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y110_SLICE_X154Y110_AQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y112_SLICE_X153Y112_BQ),
.I5(CLBLM_L_X98Y110_SLICE_X154Y110_A5Q),
.O5(CLBLM_L_X98Y110_SLICE_X154Y110_BO5),
.O6(CLBLM_L_X98Y110_SLICE_X154Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y110_SLICE_X154Y110_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y112_SLICE_X153Y112_BQ),
.I2(CLBLM_L_X98Y110_SLICE_X154Y110_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X154Y110_AO5),
.O6(CLBLM_L_X98Y110_SLICE_X154Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y110_SLICE_X155Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X155Y110_DO5),
.O6(CLBLM_L_X98Y110_SLICE_X155Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y110_SLICE_X155Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X155Y110_CO5),
.O6(CLBLM_L_X98Y110_SLICE_X155Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y110_SLICE_X155Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X155Y110_BO5),
.O6(CLBLM_L_X98Y110_SLICE_X155Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y110_SLICE_X155Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y110_SLICE_X155Y110_AO5),
.O6(CLBLM_L_X98Y110_SLICE_X155Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X154Y111_AO5),
.Q(CLBLM_L_X98Y111_SLICE_X154Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X154Y111_BO5),
.Q(CLBLM_L_X98Y111_SLICE_X154Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X154Y111_AO6),
.Q(CLBLM_L_X98Y111_SLICE_X154Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X154Y111_BO6),
.Q(CLBLM_L_X98Y111_SLICE_X154Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y111_SLICE_X154Y111_DO5),
.O6(CLBLM_L_X98Y111_SLICE_X154Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y111_SLICE_X154Y111_AQ),
.I2(CLBLM_R_X97Y112_SLICE_X152Y112_AQ),
.I3(CLBLM_L_X98Y111_SLICE_X154Y111_BQ),
.I4(CLBLM_L_X98Y111_SLICE_X154Y111_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X98Y111_SLICE_X154Y111_CO5),
.O6(CLBLM_L_X98Y111_SLICE_X154Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y111_SLICE_X154Y111_BQ),
.I2(CLBLM_L_X98Y111_SLICE_X154Y111_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y111_SLICE_X154Y111_BO5),
.O6(CLBLM_L_X98Y111_SLICE_X154Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_L_X98Y111_SLICE_X154Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y110_SLICE_X154Y110_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X97Y112_SLICE_X152Y112_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y111_SLICE_X154Y111_AO5),
.O6(CLBLM_L_X98Y111_SLICE_X154Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X155Y111_AO5),
.Q(CLBLM_L_X98Y111_SLICE_X155Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X155Y111_BO5),
.Q(CLBLM_L_X98Y111_SLICE_X155Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X155Y111_CO5),
.Q(CLBLM_L_X98Y111_SLICE_X155Y111_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X155Y111_AO6),
.Q(CLBLM_L_X98Y111_SLICE_X155Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X155Y111_BO6),
.Q(CLBLM_L_X98Y111_SLICE_X155Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y111_SLICE_X155Y111_CO6),
.Q(CLBLM_L_X98Y111_SLICE_X155Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_DLUT (
.I0(CLBLM_L_X98Y111_SLICE_X155Y111_C5Q),
.I1(CLBLM_L_X98Y111_SLICE_X155Y111_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y111_SLICE_X155Y111_BQ),
.I4(1'b1),
.I5(CLBLM_R_X95Y111_SLICE_X150Y111_AQ),
.O5(CLBLM_L_X98Y111_SLICE_X155Y111_DO5),
.O6(CLBLM_L_X98Y111_SLICE_X155Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y111_SLICE_X155Y111_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y111_SLICE_X155Y111_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y111_SLICE_X155Y111_CO5),
.O6(CLBLM_L_X98Y111_SLICE_X155Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y111_SLICE_X150Y111_AQ),
.I2(CLBLM_R_X97Y111_SLICE_X152Y111_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y111_SLICE_X155Y111_BO5),
.O6(CLBLM_L_X98Y111_SLICE_X155Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222aa0000aa)
  ) CLBLM_L_X98Y111_SLICE_X155Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y111_SLICE_X156Y111_CO6),
.I2(1'b1),
.I3(CLBLM_L_X98Y111_SLICE_X155Y111_B5Q),
.I4(CLBLL_L_X100Y111_SLICE_X157Y111_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y111_SLICE_X155Y111_AO5),
.O6(CLBLM_L_X98Y111_SLICE_X155Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y112_SLICE_X154Y112_AO5),
.Q(CLBLM_L_X98Y112_SLICE_X154Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y112_SLICE_X154Y112_BO5),
.Q(CLBLM_L_X98Y112_SLICE_X154Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y112_SLICE_X154Y112_AO6),
.Q(CLBLM_L_X98Y112_SLICE_X154Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y112_SLICE_X154Y112_BO6),
.Q(CLBLM_L_X98Y112_SLICE_X154Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X154Y112_DO5),
.O6(CLBLM_L_X98Y112_SLICE_X154Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03f3afaf03f3a0a0)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_CLUT (
.I0(CLBLL_L_X100Y112_SLICE_X156Y112_CO6),
.I1(CLBLL_L_X100Y112_SLICE_X157Y112_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y112_SLICE_X154Y112_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X97Y113_SLICE_X152Y113_BO6),
.O5(CLBLM_L_X98Y112_SLICE_X154Y112_CO5),
.O6(CLBLM_L_X98Y112_SLICE_X154Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaa00aa00a)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y112_SLICE_X155Y112_A5Q),
.I3(CLBLM_R_X97Y112_SLICE_X152Y112_B5Q),
.I4(CLBLM_L_X98Y112_SLICE_X154Y112_CO6),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X154Y112_BO5),
.O6(CLBLM_L_X98Y112_SLICE_X154Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X98Y112_SLICE_X154Y112_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y112_SLICE_X154Y112_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X100Y111_SLICE_X156Y111_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X154Y112_AO5),
.O6(CLBLM_L_X98Y112_SLICE_X154Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y112_SLICE_X155Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y112_SLICE_X155Y112_AO5),
.Q(CLBLM_L_X98Y112_SLICE_X155Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y112_SLICE_X155Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y112_SLICE_X155Y112_AO6),
.Q(CLBLM_L_X98Y112_SLICE_X155Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y112_SLICE_X155Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X155Y112_DO5),
.O6(CLBLM_L_X98Y112_SLICE_X155Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y112_SLICE_X155Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X155Y112_CO5),
.O6(CLBLM_L_X98Y112_SLICE_X155Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y112_SLICE_X155Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X155Y112_BO5),
.O6(CLBLM_L_X98Y112_SLICE_X155Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLM_L_X98Y112_SLICE_X155Y112_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y112_SLICE_X156Y112_BO6),
.I2(CLBLM_L_X98Y111_SLICE_X155Y111_C5Q),
.I3(CLBLM_L_X98Y111_SLICE_X155Y111_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y112_SLICE_X155Y112_AO5),
.O6(CLBLM_L_X98Y112_SLICE_X155Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y113_SLICE_X154Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y113_SLICE_X154Y113_AO5),
.Q(CLBLM_L_X98Y113_SLICE_X154Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y113_SLICE_X154Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y113_SLICE_X154Y113_AO6),
.Q(CLBLM_L_X98Y113_SLICE_X154Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y113_SLICE_X154Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y113_SLICE_X154Y113_DO5),
.O6(CLBLM_L_X98Y113_SLICE_X154Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5353fff053530f00)
  ) CLBLM_L_X98Y113_SLICE_X154Y113_CLUT (
.I0(CLBLM_L_X98Y115_SLICE_X154Y115_AQ),
.I1(CLBLL_L_X100Y113_SLICE_X157Y113_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y113_SLICE_X151Y113_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y114_SLICE_X154Y114_DO6),
.O5(CLBLM_L_X98Y113_SLICE_X154Y113_CO5),
.O6(CLBLM_L_X98Y113_SLICE_X154Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03aff3af03a0f3a0)
  ) CLBLM_L_X98Y113_SLICE_X154Y113_BLUT (
.I0(CLBLL_L_X100Y113_SLICE_X156Y113_DO6),
.I1(CLBLL_L_X100Y113_SLICE_X156Y113_C5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X98Y112_SLICE_X154Y112_AQ),
.I5(CLBLM_R_X95Y116_SLICE_X150Y116_CO6),
.O5(CLBLM_L_X98Y113_SLICE_X154Y113_BO5),
.O6(CLBLM_L_X98Y113_SLICE_X154Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa88882222)
  ) CLBLM_L_X98Y113_SLICE_X154Y113_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y113_SLICE_X152Y113_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y113_SLICE_X154Y113_BO6),
.I4(CLBLM_L_X98Y112_SLICE_X154Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y113_SLICE_X154Y113_AO5),
.O6(CLBLM_L_X98Y113_SLICE_X154Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y113_SLICE_X155Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y113_SLICE_X155Y113_DO5),
.O6(CLBLM_L_X98Y113_SLICE_X155Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y113_SLICE_X155Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y113_SLICE_X155Y113_CO5),
.O6(CLBLM_L_X98Y113_SLICE_X155Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y113_SLICE_X155Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y113_SLICE_X155Y113_BO5),
.O6(CLBLM_L_X98Y113_SLICE_X155Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y113_SLICE_X155Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y113_SLICE_X155Y113_AO5),
.O6(CLBLM_L_X98Y113_SLICE_X155Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y114_SLICE_X154Y114_AO5),
.Q(CLBLM_L_X98Y114_SLICE_X154Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y114_SLICE_X154Y114_BO5),
.Q(CLBLM_L_X98Y114_SLICE_X154Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y114_SLICE_X154Y114_CO5),
.Q(CLBLM_L_X98Y114_SLICE_X154Y114_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y114_SLICE_X154Y114_AO6),
.Q(CLBLM_L_X98Y114_SLICE_X154Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y114_SLICE_X154Y114_BO6),
.Q(CLBLM_L_X98Y114_SLICE_X154Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y114_SLICE_X154Y114_CO6),
.Q(CLBLM_L_X98Y114_SLICE_X154Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_DLUT (
.I0(CLBLM_L_X98Y114_SLICE_X154Y114_C5Q),
.I1(CLBLM_L_X98Y114_SLICE_X154Y114_CQ),
.I2(CLBLM_R_X97Y115_SLICE_X153Y115_AQ),
.I3(CLBLM_L_X98Y114_SLICE_X154Y114_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X154Y114_DO5),
.O6(CLBLM_L_X98Y114_SLICE_X154Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y114_SLICE_X154Y114_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y114_SLICE_X154Y114_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X154Y114_CO5),
.O6(CLBLM_L_X98Y114_SLICE_X154Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y115_SLICE_X154Y115_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X97Y115_SLICE_X153Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X154Y114_BO5),
.O6(CLBLM_L_X98Y114_SLICE_X154Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_L_X98Y114_SLICE_X154Y114_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y113_SLICE_X154Y113_A5Q),
.I2(CLBLM_R_X95Y115_SLICE_X150Y115_A5Q),
.I3(CLBLL_L_X100Y114_SLICE_X156Y114_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X154Y114_AO5),
.O6(CLBLM_L_X98Y114_SLICE_X154Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y114_SLICE_X155Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X155Y114_DO5),
.O6(CLBLM_L_X98Y114_SLICE_X155Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y114_SLICE_X155Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X155Y114_CO5),
.O6(CLBLM_L_X98Y114_SLICE_X155Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y114_SLICE_X155Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X155Y114_BO5),
.O6(CLBLM_L_X98Y114_SLICE_X155Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y114_SLICE_X155Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y114_SLICE_X155Y114_AO5),
.O6(CLBLM_L_X98Y114_SLICE_X155Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X154Y115_AO5),
.Q(CLBLM_L_X98Y115_SLICE_X154Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X154Y115_BO5),
.Q(CLBLM_L_X98Y115_SLICE_X154Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X154Y115_AO6),
.Q(CLBLM_L_X98Y115_SLICE_X154Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X154Y115_BO6),
.Q(CLBLM_L_X98Y115_SLICE_X154Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y116_SLICE_X152Y116_AQ),
.I3(CLBLM_L_X98Y115_SLICE_X154Y115_BQ),
.I4(CLBLM_L_X98Y115_SLICE_X154Y115_B5Q),
.I5(CLBLM_L_X98Y114_SLICE_X154Y114_B5Q),
.O5(CLBLM_L_X98Y115_SLICE_X154Y115_DO5),
.O6(CLBLM_L_X98Y115_SLICE_X154Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32ba109876fe54dc)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X95Y115_SLICE_X150Y115_DO6),
.I3(CLBLM_L_X98Y115_SLICE_X154Y115_A5Q),
.I4(CLBLM_L_X98Y115_SLICE_X154Y115_DO6),
.I5(CLBLL_L_X100Y115_SLICE_X156Y115_B5Q),
.O5(CLBLM_L_X98Y115_SLICE_X154Y115_CO5),
.O6(CLBLM_L_X98Y115_SLICE_X154Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y115_SLICE_X154Y115_BQ),
.I2(CLBLM_R_X97Y116_SLICE_X152Y116_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y115_SLICE_X154Y115_BO5),
.O6(CLBLM_L_X98Y115_SLICE_X154Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X98Y115_SLICE_X154Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y115_SLICE_X155Y115_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y115_SLICE_X154Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y115_SLICE_X154Y115_AO5),
.O6(CLBLM_L_X98Y115_SLICE_X154Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X155Y115_AO5),
.Q(CLBLM_L_X98Y115_SLICE_X155Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X155Y115_BO5),
.Q(CLBLM_L_X98Y115_SLICE_X155Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X155Y115_CO5),
.Q(CLBLM_L_X98Y115_SLICE_X155Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X155Y115_AO6),
.Q(CLBLM_L_X98Y115_SLICE_X155Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X155Y115_BO6),
.Q(CLBLM_L_X98Y115_SLICE_X155Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y115_SLICE_X155Y115_CO6),
.Q(CLBLM_L_X98Y115_SLICE_X155Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y115_SLICE_X155Y115_BQ),
.I3(CLBLM_L_X98Y115_SLICE_X155Y115_A5Q),
.I4(CLBLM_L_X98Y115_SLICE_X155Y115_B5Q),
.I5(CLBLM_L_X98Y114_SLICE_X154Y114_AQ),
.O5(CLBLM_L_X98Y115_SLICE_X155Y115_DO5),
.O6(CLBLM_L_X98Y115_SLICE_X155Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f0f00000)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_CLUT (
.I0(CLBLM_L_X98Y115_SLICE_X155Y115_C5Q),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y115_SLICE_X143Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y115_SLICE_X155Y115_CO5),
.O6(CLBLM_L_X98Y115_SLICE_X155Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y115_SLICE_X155Y115_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y114_SLICE_X154Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y115_SLICE_X155Y115_BO5),
.O6(CLBLM_L_X98Y115_SLICE_X155Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X98Y115_SLICE_X155Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y115_SLICE_X152Y115_AQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y115_SLICE_X155Y115_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y115_SLICE_X155Y115_AO5),
.O6(CLBLM_L_X98Y115_SLICE_X155Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y116_SLICE_X154Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y116_SLICE_X154Y116_DO5),
.O6(CLBLM_L_X98Y116_SLICE_X154Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y116_SLICE_X154Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y116_SLICE_X154Y116_CO5),
.O6(CLBLM_L_X98Y116_SLICE_X154Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y116_SLICE_X154Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y116_SLICE_X154Y116_BO5),
.O6(CLBLM_L_X98Y116_SLICE_X154Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00acf0ac0facffac)
  ) CLBLM_L_X98Y116_SLICE_X154Y116_ALUT (
.I0(CLBLL_L_X100Y116_SLICE_X157Y116_DO6),
.I1(CLBLM_R_X93Y116_SLICE_X146Y116_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X100Y114_SLICE_X156Y114_AQ),
.I5(CLBLL_L_X100Y116_SLICE_X157Y116_B5Q),
.O5(CLBLM_L_X98Y116_SLICE_X154Y116_AO5),
.O6(CLBLM_L_X98Y116_SLICE_X154Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y116_SLICE_X155Y116_AO5),
.Q(CLBLM_L_X98Y116_SLICE_X155Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y116_SLICE_X155Y116_BO5),
.Q(CLBLM_L_X98Y116_SLICE_X155Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y116_SLICE_X155Y116_AO6),
.Q(CLBLM_L_X98Y116_SLICE_X155Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y116_SLICE_X155Y116_BO6),
.Q(CLBLM_L_X98Y116_SLICE_X155Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y116_SLICE_X153Y116_B5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y116_SLICE_X155Y116_BQ),
.I4(CLBLM_L_X98Y116_SLICE_X155Y116_B5Q),
.I5(CLBLL_L_X100Y117_SLICE_X156Y117_A5Q),
.O5(CLBLM_L_X98Y116_SLICE_X155Y116_DO5),
.O6(CLBLM_L_X98Y116_SLICE_X155Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777444430fc30fc)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_CLUT (
.I0(CLBLM_L_X98Y115_SLICE_X155Y115_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X92Y116_SLICE_X144Y116_DO6),
.I3(CLBLM_L_X98Y116_SLICE_X155Y116_A5Q),
.I4(CLBLM_L_X98Y116_SLICE_X155Y116_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X98Y116_SLICE_X155Y116_CO5),
.O6(CLBLM_L_X98Y116_SLICE_X155Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y116_SLICE_X155Y116_BQ),
.I2(1'b1),
.I3(CLBLL_L_X100Y117_SLICE_X156Y117_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y116_SLICE_X155Y116_BO5),
.O6(CLBLM_L_X98Y116_SLICE_X155Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaa00aa00a)
  ) CLBLM_L_X98Y116_SLICE_X155Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X92Y116_SLICE_X145Y116_A5Q),
.I3(CLBLM_R_X97Y116_SLICE_X153Y116_B5Q),
.I4(CLBLL_L_X100Y116_SLICE_X156Y116_CO6),
.I5(1'b1),
.O5(CLBLM_L_X98Y116_SLICE_X155Y116_AO5),
.O6(CLBLM_L_X98Y116_SLICE_X155Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y117_SLICE_X154Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y117_SLICE_X154Y117_DO5),
.O6(CLBLM_L_X98Y117_SLICE_X154Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y117_SLICE_X154Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y117_SLICE_X154Y117_CO5),
.O6(CLBLM_L_X98Y117_SLICE_X154Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y117_SLICE_X154Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y117_SLICE_X154Y117_BO5),
.O6(CLBLM_L_X98Y117_SLICE_X154Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f90609f9f60906)
  ) CLBLM_L_X98Y117_SLICE_X154Y117_ALUT (
.I0(CLBLM_R_X97Y117_SLICE_X153Y117_BQ),
.I1(CLBLM_R_X97Y118_SLICE_X153Y118_BQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y117_SLICE_X153Y117_C5Q),
.I4(CLBLL_L_X100Y118_SLICE_X157Y118_C5Q),
.I5(CLBLM_R_X97Y117_SLICE_X152Y117_B5Q),
.O5(CLBLM_L_X98Y117_SLICE_X154Y117_AO5),
.O6(CLBLM_L_X98Y117_SLICE_X154Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y117_SLICE_X155Y117_AO5),
.Q(CLBLM_L_X98Y117_SLICE_X155Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y117_SLICE_X155Y117_BO5),
.Q(CLBLM_L_X98Y117_SLICE_X155Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y117_SLICE_X155Y117_AO6),
.Q(CLBLM_L_X98Y117_SLICE_X155Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y117_SLICE_X155Y117_BO6),
.Q(CLBLM_L_X98Y117_SLICE_X155Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_DLUT (
.I0(CLBLM_L_X94Y116_SLICE_X149Y116_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y119_SLICE_X155Y119_B5Q),
.I3(CLBLM_L_X98Y117_SLICE_X155Y117_BQ),
.I4(CLBLM_L_X98Y117_SLICE_X155Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y117_SLICE_X155Y117_DO5),
.O6(CLBLM_L_X98Y117_SLICE_X155Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033aaf0ff33aaf0)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_CLUT (
.I0(CLBLM_L_X98Y117_SLICE_X155Y117_DO6),
.I1(CLBLL_L_X100Y118_SLICE_X157Y118_A5Q),
.I2(CLBLM_R_X93Y117_SLICE_X146Y117_CO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y117_SLICE_X155Y117_AQ),
.O5(CLBLM_L_X98Y117_SLICE_X155Y117_CO5),
.O6(CLBLM_L_X98Y117_SLICE_X155Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y117_SLICE_X155Y117_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X94Y116_SLICE_X149Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y117_SLICE_X155Y117_BO5),
.O6(CLBLM_L_X98Y117_SLICE_X155Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa000a0a0a0a)
  ) CLBLM_L_X98Y117_SLICE_X155Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y117_SLICE_X155Y117_AQ),
.I3(CLBLL_L_X100Y114_SLICE_X156Y114_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y117_SLICE_X155Y117_AO5),
.O6(CLBLM_L_X98Y117_SLICE_X155Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X154Y119_AO5),
.Q(CLBLM_L_X98Y119_SLICE_X154Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X154Y119_CO5),
.Q(CLBLM_L_X98Y119_SLICE_X154Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X154Y119_AO6),
.Q(CLBLM_L_X98Y119_SLICE_X154Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X154Y119_BO6),
.Q(CLBLM_L_X98Y119_SLICE_X154Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12ed21ed21de12)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_DLUT (
.I0(CLBLM_L_X98Y120_SLICE_X154Y120_CQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X97Y118_SLICE_X153Y118_C5Q),
.I3(CLBLL_L_X100Y118_SLICE_X157Y118_BQ),
.I4(CLBLM_L_X98Y119_SLICE_X154Y119_BQ),
.I5(CLBLM_L_X98Y119_SLICE_X154Y119_B5Q),
.O5(CLBLM_L_X98Y119_SLICE_X154Y119_DO5),
.O6(CLBLM_L_X98Y119_SLICE_X154Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696f000f000)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_CLUT (
.I0(CLBLM_L_X98Y120_SLICE_X154Y120_CQ),
.I1(CLBLM_L_X98Y119_SLICE_X154Y119_B5Q),
.I2(CLBLM_R_X97Y118_SLICE_X153Y118_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y119_SLICE_X154Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y119_SLICE_X154Y119_CO5),
.O6(CLBLM_L_X98Y119_SLICE_X154Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha088aa88a0880088)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y118_SLICE_X142Y118_CO6),
.I2(CLBLM_L_X98Y119_SLICE_X154Y119_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y119_SLICE_X154Y119_CO6),
.O5(CLBLM_L_X98Y119_SLICE_X154Y119_BO5),
.O6(CLBLM_L_X98Y119_SLICE_X154Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X98Y119_SLICE_X154Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y119_SLICE_X154Y119_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X97Y122_SLICE_X152Y122_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y119_SLICE_X154Y119_AO5),
.O6(CLBLM_L_X98Y119_SLICE_X154Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X155Y119_BO5),
.Q(CLBLM_L_X98Y119_SLICE_X155Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X155Y119_CO5),
.Q(CLBLM_L_X98Y119_SLICE_X155Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X155Y119_AO6),
.Q(CLBLM_L_X98Y119_SLICE_X155Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X155Y119_BO6),
.Q(CLBLM_L_X98Y119_SLICE_X155Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y119_SLICE_X155Y119_CO6),
.Q(CLBLM_L_X98Y119_SLICE_X155Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_DLUT (
.I0(CLBLM_L_X98Y119_SLICE_X155Y119_C5Q),
.I1(CLBLM_L_X98Y119_SLICE_X155Y119_CQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y120_SLICE_X155Y120_A5Q),
.I4(CLBLM_R_X97Y119_SLICE_X152Y119_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X98Y119_SLICE_X155Y119_DO5),
.O6(CLBLM_L_X98Y119_SLICE_X155Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y119_SLICE_X155Y119_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y119_SLICE_X152Y119_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y119_SLICE_X155Y119_CO5),
.O6(CLBLM_L_X98Y119_SLICE_X155Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y119_SLICE_X155Y119_AQ),
.I3(1'b1),
.I4(CLBLM_L_X98Y117_SLICE_X155Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y119_SLICE_X155Y119_BO5),
.O6(CLBLM_L_X98Y119_SLICE_X155Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a28080aa228800)
  ) CLBLM_L_X98Y119_SLICE_X155Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y119_SLICE_X154Y119_A5Q),
.I3(CLBLL_L_X100Y119_SLICE_X156Y119_AO6),
.I4(CLBLM_L_X92Y118_SLICE_X144Y118_BO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y119_SLICE_X155Y119_AO5),
.O6(CLBLM_L_X98Y119_SLICE_X155Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X154Y120_BO5),
.Q(CLBLM_L_X98Y120_SLICE_X154Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X154Y120_CO5),
.Q(CLBLM_L_X98Y120_SLICE_X154Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X154Y120_AO6),
.Q(CLBLM_L_X98Y120_SLICE_X154Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X154Y120_CO6),
.Q(CLBLM_L_X98Y120_SLICE_X154Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3276bafe105498dc)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y125_SLICE_X163Y125_DO6),
.I3(CLBLM_R_X97Y120_SLICE_X153Y120_B5Q),
.I4(CLBLL_L_X100Y122_SLICE_X157Y122_B5Q),
.I5(CLBLM_L_X98Y119_SLICE_X155Y119_DO6),
.O5(CLBLM_L_X98Y120_SLICE_X154Y120_DO5),
.O6(CLBLM_L_X98Y120_SLICE_X154Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f000f000)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_CLUT (
.I0(CLBLM_L_X98Y119_SLICE_X154Y119_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y121_SLICE_X154Y121_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y120_SLICE_X154Y120_CO5),
.O6(CLBLM_L_X98Y120_SLICE_X154Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y120_SLICE_X154Y120_A5Q),
.I2(CLBLM_L_X98Y120_SLICE_X154Y120_AQ),
.I3(CLBLM_L_X98Y121_SLICE_X154Y121_DQ),
.I4(CLBLM_L_X98Y120_SLICE_X154Y120_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y120_SLICE_X154Y120_BO5),
.O6(CLBLM_L_X98Y120_SLICE_X154Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a8080aa0aa000)
  ) CLBLM_L_X98Y120_SLICE_X154Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y122_SLICE_X152Y122_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y120_SLICE_X154Y120_BO6),
.I4(CLBLM_R_X89Y120_SLICE_X140Y120_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y120_SLICE_X154Y120_AO5),
.O6(CLBLM_L_X98Y120_SLICE_X154Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X155Y120_AO5),
.Q(CLBLM_L_X98Y120_SLICE_X155Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X155Y120_BO5),
.Q(CLBLM_L_X98Y120_SLICE_X155Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X155Y120_AO6),
.Q(CLBLM_L_X98Y120_SLICE_X155Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y120_SLICE_X155Y120_BO6),
.Q(CLBLM_L_X98Y120_SLICE_X155Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_DLUT (
.I0(CLBLM_L_X98Y120_SLICE_X155Y120_BQ),
.I1(CLBLM_L_X98Y120_SLICE_X155Y120_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y118_SLICE_X158Y118_A5Q),
.I4(CLBLM_L_X98Y120_SLICE_X155Y120_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y120_SLICE_X155Y120_DO5),
.O6(CLBLM_L_X98Y120_SLICE_X155Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_CLUT (
.I0(CLBLM_L_X98Y120_SLICE_X154Y120_AQ),
.I1(CLBLM_L_X98Y121_SLICE_X154Y121_DQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X101Y119_SLICE_X158Y119_CQ),
.I4(CLBLM_L_X98Y120_SLICE_X154Y120_C5Q),
.I5(CLBLM_L_X98Y120_SLICE_X154Y120_A5Q),
.O5(CLBLM_L_X98Y120_SLICE_X155Y120_CO5),
.O6(CLBLM_L_X98Y120_SLICE_X155Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y120_SLICE_X155Y120_BQ),
.I2(CLBLM_L_X98Y120_SLICE_X155Y120_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y120_SLICE_X155Y120_BO5),
.O6(CLBLM_L_X98Y120_SLICE_X155Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y120_SLICE_X155Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y118_SLICE_X158Y118_A5Q),
.I2(CLBLM_L_X98Y119_SLICE_X155Y119_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y120_SLICE_X155Y120_AO5),
.O6(CLBLM_L_X98Y120_SLICE_X155Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X154Y121_AO5),
.Q(CLBLM_L_X98Y121_SLICE_X154Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X154Y121_DO5),
.Q(CLBLM_L_X98Y121_SLICE_X154Y121_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X154Y121_AO6),
.Q(CLBLM_L_X98Y121_SLICE_X154Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X154Y121_BO5),
.Q(CLBLM_L_X98Y121_SLICE_X154Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X154Y121_CO6),
.Q(CLBLM_L_X98Y121_SLICE_X154Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X154Y121_DO6),
.Q(CLBLM_L_X98Y121_SLICE_X154Y121_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0c0c0c0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_DLUT (
.I0(CLBLM_L_X98Y120_SLICE_X154Y120_AQ),
.I1(CLBLM_L_X98Y122_SLICE_X154Y122_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y121_SLICE_X154Y121_DO5),
.O6(CLBLM_L_X98Y121_SLICE_X154Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0f080c0b0308000)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_CLUT (
.I0(CLBLM_L_X98Y121_SLICE_X154Y121_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X93Y122_SLICE_X147Y122_DO6),
.I5(CLBLM_L_X98Y121_SLICE_X155Y121_AO6),
.O5(CLBLM_L_X98Y121_SLICE_X154Y121_CO5),
.O6(CLBLM_L_X98Y121_SLICE_X154Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33ca0a0a0a0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y121_SLICE_X154Y121_BQ),
.I2(CLBLM_L_X98Y121_SLICE_X154Y121_D5Q),
.I3(CLBLM_L_X98Y122_SLICE_X154Y122_BQ),
.I4(CLBLM_R_X97Y122_SLICE_X152Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y121_SLICE_X154Y121_BO5),
.O6(CLBLM_L_X98Y121_SLICE_X154Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y121_SLICE_X154Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y121_SLICE_X154Y121_A5Q),
.I2(CLBLL_L_X100Y121_SLICE_X156Y121_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y121_SLICE_X154Y121_AO5),
.O6(CLBLM_L_X98Y121_SLICE_X154Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X155Y121_BO5),
.Q(CLBLM_L_X98Y121_SLICE_X155Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X155Y121_CO5),
.Q(CLBLM_L_X98Y121_SLICE_X155Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X155Y121_AO5),
.Q(CLBLM_L_X98Y121_SLICE_X155Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X155Y121_BO6),
.Q(CLBLM_L_X98Y121_SLICE_X155Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y121_SLICE_X155Y121_CO6),
.Q(CLBLM_L_X98Y121_SLICE_X155Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_DLUT (
.I0(CLBLL_L_X102Y120_SLICE_X160Y120_D5Q),
.I1(CLBLM_L_X98Y121_SLICE_X155Y121_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y121_SLICE_X154Y121_CQ),
.I4(CLBLM_L_X98Y121_SLICE_X155Y121_B5Q),
.I5(CLBLM_L_X98Y121_SLICE_X155Y121_AQ),
.O5(CLBLM_L_X98Y121_SLICE_X155Y121_DO5),
.O6(CLBLM_L_X98Y121_SLICE_X155Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f0f00000)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_CLUT (
.I0(CLBLM_L_X98Y121_SLICE_X154Y121_CQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y121_SLICE_X157Y121_CQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y121_SLICE_X155Y121_CO5),
.O6(CLBLM_L_X98Y121_SLICE_X155Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y121_SLICE_X155Y121_CQ),
.I3(1'b1),
.I4(CLBLM_L_X98Y123_SLICE_X155Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y121_SLICE_X155Y121_BO5),
.O6(CLBLM_L_X98Y121_SLICE_X155Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c88888888)
  ) CLBLM_L_X98Y121_SLICE_X155Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y121_SLICE_X155Y121_B5Q),
.I2(CLBLM_L_X98Y121_SLICE_X155Y121_CQ),
.I3(CLBLM_L_X98Y121_SLICE_X155Y121_AQ),
.I4(CLBLM_L_X98Y121_SLICE_X154Y121_CQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y121_SLICE_X155Y121_AO5),
.O6(CLBLM_L_X98Y121_SLICE_X155Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X154Y122_AO5),
.Q(CLBLM_L_X98Y122_SLICE_X154Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X154Y122_BO5),
.Q(CLBLM_L_X98Y122_SLICE_X154Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X154Y122_AO6),
.Q(CLBLM_L_X98Y122_SLICE_X154Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X154Y122_BO6),
.Q(CLBLM_L_X98Y122_SLICE_X154Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X97Y122_SLICE_X153Y122_AQ),
.I2(CLBLM_R_X101Y123_SLICE_X159Y123_CQ),
.I3(CLBLM_L_X98Y123_SLICE_X154Y123_CQ),
.I4(CLBLM_L_X98Y122_SLICE_X154Y122_B5Q),
.I5(CLBLM_R_X97Y122_SLICE_X152Y122_CQ),
.O5(CLBLM_L_X98Y122_SLICE_X154Y122_DO5),
.O6(CLBLM_L_X98Y122_SLICE_X154Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_CLUT (
.I0(CLBLM_R_X97Y122_SLICE_X152Y122_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X98Y122_SLICE_X154Y122_BQ),
.I3(CLBLM_L_X98Y121_SLICE_X154Y121_D5Q),
.I4(CLBLM_R_X101Y123_SLICE_X159Y123_C5Q),
.I5(CLBLM_L_X98Y121_SLICE_X154Y121_BQ),
.O5(CLBLM_L_X98Y122_SLICE_X154Y122_CO5),
.O6(CLBLM_L_X98Y122_SLICE_X154Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y123_SLICE_X154Y123_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X97Y122_SLICE_X152Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y122_SLICE_X154Y122_BO5),
.O6(CLBLM_L_X98Y122_SLICE_X154Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y122_SLICE_X154Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y122_SLICE_X154Y122_A5Q),
.I2(CLBLM_L_X98Y121_SLICE_X154Y121_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y122_SLICE_X154Y122_AO5),
.O6(CLBLM_L_X98Y122_SLICE_X154Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X155Y122_AO5),
.Q(CLBLM_L_X98Y122_SLICE_X155Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X155Y122_BO5),
.Q(CLBLM_L_X98Y122_SLICE_X155Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X155Y122_AO6),
.Q(CLBLM_L_X98Y122_SLICE_X155Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y122_SLICE_X155Y122_BO6),
.Q(CLBLM_L_X98Y122_SLICE_X155Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_DLUT (
.I0(CLBLM_L_X98Y122_SLICE_X155Y122_BQ),
.I1(CLBLM_R_X97Y122_SLICE_X153Y122_B5Q),
.I2(CLBLL_L_X100Y123_SLICE_X156Y123_BQ),
.I3(1'b1),
.I4(CLBLM_L_X98Y122_SLICE_X155Y122_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X98Y122_SLICE_X155Y122_DO5),
.O6(CLBLM_L_X98Y122_SLICE_X155Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f50500cfc0cfc)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_CLUT (
.I0(CLBLM_L_X98Y122_SLICE_X155Y122_A5Q),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y122_SLICE_X152Y122_D5Q),
.I4(CLBLM_L_X98Y122_SLICE_X155Y122_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X98Y122_SLICE_X155Y122_CO5),
.O6(CLBLM_L_X98Y122_SLICE_X155Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y122_SLICE_X155Y122_BQ),
.I2(1'b1),
.I3(CLBLL_L_X100Y123_SLICE_X156Y123_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y122_SLICE_X155Y122_BO5),
.O6(CLBLM_L_X98Y122_SLICE_X155Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y122_SLICE_X155Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y122_SLICE_X155Y122_A5Q),
.I2(CLBLM_R_X97Y124_SLICE_X152Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y122_SLICE_X155Y122_AO5),
.O6(CLBLM_L_X98Y122_SLICE_X155Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X154Y123_BO5),
.Q(CLBLM_L_X98Y123_SLICE_X154Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X154Y123_CO5),
.Q(CLBLM_L_X98Y123_SLICE_X154Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X154Y123_AO6),
.Q(CLBLM_L_X98Y123_SLICE_X154Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X154Y123_CO6),
.Q(CLBLM_L_X98Y123_SLICE_X154Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_DLUT (
.I0(CLBLM_L_X98Y123_SLICE_X154Y123_C5Q),
.I1(CLBLM_L_X98Y123_SLICE_X154Y123_AQ),
.I2(CLBLL_L_X102Y124_SLICE_X160Y124_D5Q),
.I3(CLBLM_L_X98Y123_SLICE_X155Y123_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y123_SLICE_X154Y123_A5Q),
.O5(CLBLM_L_X98Y123_SLICE_X154Y123_DO5),
.O6(CLBLM_L_X98Y123_SLICE_X154Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000a0a0a0a0)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_CLUT (
.I0(CLBLM_L_X98Y123_SLICE_X155Y123_CQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y122_SLICE_X152Y122_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y123_SLICE_X154Y123_CO5),
.O6(CLBLM_L_X98Y123_SLICE_X154Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y123_SLICE_X155Y123_CQ),
.I2(CLBLM_L_X98Y123_SLICE_X154Y123_AQ),
.I3(CLBLM_L_X98Y123_SLICE_X154Y123_A5Q),
.I4(CLBLM_L_X98Y123_SLICE_X154Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y123_SLICE_X154Y123_BO5),
.O6(CLBLM_L_X98Y123_SLICE_X154Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa8a2a0aa0802000)
  ) CLBLM_L_X98Y123_SLICE_X154Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y123_SLICE_X154Y123_BO6),
.I4(CLBLM_L_X98Y122_SLICE_X154Y122_A5Q),
.I5(CLBLM_R_X93Y123_SLICE_X146Y123_DO6),
.O5(CLBLM_L_X98Y123_SLICE_X154Y123_AO5),
.O6(CLBLM_L_X98Y123_SLICE_X154Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X155Y123_BO5),
.Q(CLBLM_L_X98Y123_SLICE_X155Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X155Y123_CO5),
.Q(CLBLM_L_X98Y123_SLICE_X155Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X155Y123_AO6),
.Q(CLBLM_L_X98Y123_SLICE_X155Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y123_SLICE_X155Y123_CO6),
.Q(CLBLM_L_X98Y123_SLICE_X155Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_DLUT (
.I0(CLBLM_L_X98Y123_SLICE_X155Y123_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y124_SLICE_X160Y124_DQ),
.I3(CLBLM_L_X98Y123_SLICE_X155Y123_A5Q),
.I4(CLBLM_L_X98Y123_SLICE_X155Y123_AQ),
.I5(CLBLM_L_X98Y121_SLICE_X155Y121_BQ),
.O5(CLBLM_L_X98Y123_SLICE_X155Y123_DO5),
.O6(CLBLM_L_X98Y123_SLICE_X155Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000a0a0a0a0)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_CLUT (
.I0(CLBLM_L_X98Y121_SLICE_X155Y121_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X98Y123_SLICE_X154Y123_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y123_SLICE_X155Y123_CO5),
.O6(CLBLM_L_X98Y123_SLICE_X155Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y123_SLICE_X155Y123_A5Q),
.I2(CLBLM_L_X98Y123_SLICE_X155Y123_AQ),
.I3(CLBLM_L_X98Y121_SLICE_X155Y121_BQ),
.I4(CLBLM_L_X98Y123_SLICE_X155Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y123_SLICE_X155Y123_BO5),
.O6(CLBLM_L_X98Y123_SLICE_X155Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa8a2a0aa0802000)
  ) CLBLM_L_X98Y123_SLICE_X155Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y123_SLICE_X155Y123_BO6),
.I4(CLBLM_L_X98Y121_SLICE_X154Y121_AQ),
.I5(CLBLM_R_X93Y123_SLICE_X147Y123_DO6),
.O5(CLBLM_L_X98Y123_SLICE_X155Y123_AO5),
.O6(CLBLM_L_X98Y123_SLICE_X155Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y124_SLICE_X154Y124_AO5),
.Q(CLBLM_L_X98Y124_SLICE_X154Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y124_SLICE_X154Y124_BO5),
.Q(CLBLM_L_X98Y124_SLICE_X154Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y124_SLICE_X154Y124_AO6),
.Q(CLBLM_L_X98Y124_SLICE_X154Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y124_SLICE_X154Y124_BO6),
.Q(CLBLM_L_X98Y124_SLICE_X154Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y124_SLICE_X154Y124_BQ),
.I3(CLBLM_L_X98Y124_SLICE_X154Y124_A5Q),
.I4(CLBLM_L_X98Y124_SLICE_X154Y124_B5Q),
.I5(CLBLL_L_X100Y125_SLICE_X157Y125_CQ),
.O5(CLBLM_L_X98Y124_SLICE_X154Y124_DO5),
.O6(CLBLM_L_X98Y124_SLICE_X154Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500ffccccf0f0)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_CLUT (
.I0(CLBLL_L_X100Y123_SLICE_X157Y123_AQ),
.I1(CLBLM_R_X97Y123_SLICE_X153Y123_DO6),
.I2(CLBLL_L_X100Y125_SLICE_X156Y125_CO6),
.I3(CLBLM_R_X97Y123_SLICE_X153Y123_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y124_SLICE_X154Y124_CO5),
.O6(CLBLM_L_X98Y124_SLICE_X154Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y124_SLICE_X154Y124_BQ),
.I2(1'b1),
.I3(CLBLL_L_X100Y125_SLICE_X157Y125_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y124_SLICE_X154Y124_BO5),
.O6(CLBLM_L_X98Y124_SLICE_X154Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X98Y124_SLICE_X154Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y124_SLICE_X154Y124_B5Q),
.I2(1'b1),
.I3(CLBLL_L_X100Y124_SLICE_X157Y124_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y124_SLICE_X154Y124_AO5),
.O6(CLBLM_L_X98Y124_SLICE_X154Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y124_SLICE_X155Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y124_SLICE_X155Y124_DO5),
.O6(CLBLM_L_X98Y124_SLICE_X155Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y124_SLICE_X155Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y124_SLICE_X155Y124_CO5),
.O6(CLBLM_L_X98Y124_SLICE_X155Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y124_SLICE_X155Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y124_SLICE_X155Y124_BO5),
.O6(CLBLM_L_X98Y124_SLICE_X155Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y124_SLICE_X155Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y124_SLICE_X155Y124_AO5),
.O6(CLBLM_L_X98Y124_SLICE_X155Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_AO5),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_BO5),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_CO5),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_DO5),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_AO6),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_BO6),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_CO6),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X154Y125_DO6),
.Q(CLBLM_L_X98Y125_SLICE_X154Y125_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99990000f00f0000)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_DLUT (
.I0(CLBLM_R_X97Y126_SLICE_X153Y126_C5Q),
.I1(CLBLM_R_X95Y125_SLICE_X150Y125_B5Q),
.I2(CLBLM_L_X98Y125_SLICE_X154Y125_DQ),
.I3(CLBLM_R_X95Y124_SLICE_X151Y124_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X98Y125_SLICE_X154Y125_DO5),
.O6(CLBLM_L_X98Y125_SLICE_X154Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f090909090)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_CLUT (
.I0(CLBLL_L_X100Y124_SLICE_X157Y124_B5Q),
.I1(CLBLL_L_X100Y126_SLICE_X156Y126_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X97Y125_SLICE_X153Y125_CO6),
.I5(1'b1),
.O5(CLBLM_L_X98Y125_SLICE_X154Y125_CO5),
.O6(CLBLM_L_X98Y125_SLICE_X154Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y123_SLICE_X157Y123_AQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y125_SLICE_X154Y125_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y125_SLICE_X154Y125_BO5),
.O6(CLBLM_L_X98Y125_SLICE_X154Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa28822882)
  ) CLBLM_L_X98Y125_SLICE_X154Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y127_SLICE_X155Y127_B5Q),
.I2(CLBLM_R_X101Y126_SLICE_X159Y126_A5Q),
.I3(CLBLM_L_X98Y128_SLICE_X154Y128_A5Q),
.I4(CLBLM_R_X97Y124_SLICE_X153Y124_AO6),
.I5(1'b1),
.O5(CLBLM_L_X98Y125_SLICE_X154Y125_AO5),
.O6(CLBLM_L_X98Y125_SLICE_X154Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X155Y125_BO5),
.Q(CLBLM_L_X98Y125_SLICE_X155Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X155Y125_CO5),
.Q(CLBLM_L_X98Y125_SLICE_X155Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X155Y125_AO6),
.Q(CLBLM_L_X98Y125_SLICE_X155Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y125_SLICE_X155Y125_CO6),
.Q(CLBLM_L_X98Y125_SLICE_X155Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_DLUT (
.I0(CLBLM_L_X98Y125_SLICE_X155Y125_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X98Y125_SLICE_X155Y125_A5Q),
.I3(CLBLM_L_X98Y125_SLICE_X155Y125_AQ),
.I4(CLBLM_L_X98Y125_SLICE_X154Y125_DQ),
.I5(CLBLM_L_X98Y125_SLICE_X155Y125_CQ),
.O5(CLBLM_L_X98Y125_SLICE_X155Y125_DO5),
.O6(CLBLM_L_X98Y125_SLICE_X155Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y125_SLICE_X155Y125_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X98Y125_SLICE_X155Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y125_SLICE_X155Y125_CO5),
.O6(CLBLM_L_X98Y125_SLICE_X155Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y125_SLICE_X155Y125_A5Q),
.I2(CLBLM_L_X98Y125_SLICE_X155Y125_AQ),
.I3(CLBLM_L_X98Y125_SLICE_X155Y125_CQ),
.I4(CLBLM_L_X98Y125_SLICE_X155Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y125_SLICE_X155Y125_BO5),
.O6(CLBLM_L_X98Y125_SLICE_X155Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa8a2a0aa0802000)
  ) CLBLM_L_X98Y125_SLICE_X155Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y125_SLICE_X155Y125_BO6),
.I4(CLBLM_L_X98Y126_SLICE_X154Y126_AQ),
.I5(CLBLM_R_X103Y126_SLICE_X162Y126_DO6),
.O5(CLBLM_L_X98Y125_SLICE_X155Y125_AO5),
.O6(CLBLM_L_X98Y125_SLICE_X155Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X154Y126_AO5),
.Q(CLBLM_L_X98Y126_SLICE_X154Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X154Y126_BO5),
.Q(CLBLM_L_X98Y126_SLICE_X154Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X154Y126_AO6),
.Q(CLBLM_L_X98Y126_SLICE_X154Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X154Y126_BO6),
.Q(CLBLM_L_X98Y126_SLICE_X154Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y126_SLICE_X154Y126_DO5),
.O6(CLBLM_L_X98Y126_SLICE_X154Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055e4e4aaffe4e4)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X100Y127_SLICE_X156Y127_CO6),
.I2(CLBLM_R_X97Y125_SLICE_X153Y125_DO6),
.I3(CLBLM_R_X97Y125_SLICE_X152Y125_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y125_SLICE_X154Y125_BQ),
.O5(CLBLM_L_X98Y126_SLICE_X154Y126_CO5),
.O6(CLBLM_L_X98Y126_SLICE_X154Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y125_SLICE_X154Y125_C5Q),
.I2(1'b1),
.I3(CLBLL_L_X100Y126_SLICE_X156Y126_B5Q),
.I4(CLBLM_L_X98Y126_SLICE_X154Y126_CO6),
.I5(1'b1),
.O5(CLBLM_L_X98Y126_SLICE_X154Y126_BO5),
.O6(CLBLM_L_X98Y126_SLICE_X154Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y126_SLICE_X154Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y126_SLICE_X154Y126_A5Q),
.I2(CLBLM_R_X97Y129_SLICE_X152Y129_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y126_SLICE_X154Y126_AO5),
.O6(CLBLM_L_X98Y126_SLICE_X154Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X155Y126_BO5),
.Q(CLBLM_L_X98Y126_SLICE_X155Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X155Y126_CO5),
.Q(CLBLM_L_X98Y126_SLICE_X155Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X155Y126_AO6),
.Q(CLBLM_L_X98Y126_SLICE_X155Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y126_SLICE_X155Y126_CO6),
.Q(CLBLM_L_X98Y126_SLICE_X155Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_DLUT (
.I0(CLBLM_L_X98Y126_SLICE_X155Y126_C5Q),
.I1(CLBLM_L_X98Y126_SLICE_X155Y126_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y126_SLICE_X155Y126_A5Q),
.I4(CLBLM_L_X98Y126_SLICE_X155Y126_AQ),
.I5(CLBLM_R_X97Y126_SLICE_X153Y126_C5Q),
.O5(CLBLM_L_X98Y126_SLICE_X155Y126_DO5),
.O6(CLBLM_L_X98Y126_SLICE_X155Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y126_SLICE_X155Y126_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X98Y126_SLICE_X155Y126_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y126_SLICE_X155Y126_CO5),
.O6(CLBLM_L_X98Y126_SLICE_X155Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_BLUT (
.I0(CLBLM_L_X98Y126_SLICE_X155Y126_CQ),
.I1(CLBLM_L_X98Y126_SLICE_X155Y126_A5Q),
.I2(CLBLM_L_X98Y126_SLICE_X155Y126_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y126_SLICE_X155Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y126_SLICE_X155Y126_BO5),
.O6(CLBLM_L_X98Y126_SLICE_X155Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a28080aa228800)
  ) CLBLM_L_X98Y126_SLICE_X155Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y126_SLICE_X154Y126_A5Q),
.I3(CLBLM_L_X98Y126_SLICE_X155Y126_BO6),
.I4(CLBLL_L_X102Y127_SLICE_X161Y127_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y126_SLICE_X155Y126_AO5),
.O6(CLBLM_L_X98Y126_SLICE_X155Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X154Y127_AO5),
.Q(CLBLM_L_X98Y127_SLICE_X154Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X154Y127_BO5),
.Q(CLBLM_L_X98Y127_SLICE_X154Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X154Y127_AO6),
.Q(CLBLM_L_X98Y127_SLICE_X154Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X154Y127_BO6),
.Q(CLBLM_L_X98Y127_SLICE_X154Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bb11bbfafa5050)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y126_SLICE_X152Y126_A5Q),
.I2(CLBLL_L_X100Y127_SLICE_X157Y127_CO6),
.I3(CLBLM_L_X98Y127_SLICE_X154Y127_A5Q),
.I4(CLBLM_R_X97Y126_SLICE_X152Y126_CO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y127_SLICE_X154Y127_DO5),
.O6(CLBLM_L_X98Y127_SLICE_X154Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22227777fa50fa50)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X98Y127_SLICE_X154Y127_AQ),
.I2(CLBLM_R_X101Y129_SLICE_X158Y129_DO6),
.I3(CLBLM_R_X97Y127_SLICE_X152Y127_DO6),
.I4(CLBLM_R_X97Y127_SLICE_X153Y127_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y127_SLICE_X154Y127_CO5),
.O6(CLBLM_L_X98Y127_SLICE_X154Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y127_SLICE_X154Y127_DO6),
.I2(CLBLL_L_X100Y127_SLICE_X156Y127_A5Q),
.I3(CLBLM_L_X98Y126_SLICE_X154Y126_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y127_SLICE_X154Y127_BO5),
.O6(CLBLM_L_X98Y127_SLICE_X154Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X98Y127_SLICE_X154Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y127_SLICE_X154Y127_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y125_SLICE_X154Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y127_SLICE_X154Y127_AO5),
.O6(CLBLM_L_X98Y127_SLICE_X154Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X155Y127_AO5),
.Q(CLBLM_L_X98Y127_SLICE_X155Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X155Y127_BO5),
.Q(CLBLM_L_X98Y127_SLICE_X155Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X155Y127_AO6),
.Q(CLBLM_L_X98Y127_SLICE_X155Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y127_SLICE_X155Y127_BO6),
.Q(CLBLM_L_X98Y127_SLICE_X155Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y127_SLICE_X155Y127_DO5),
.O6(CLBLM_L_X98Y127_SLICE_X155Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X98Y128_SLICE_X154Y128_CQ),
.I2(CLBLM_L_X98Y127_SLICE_X155Y127_BQ),
.I3(CLBLM_R_X101Y128_SLICE_X158Y128_AQ),
.I4(CLBLM_L_X98Y127_SLICE_X155Y127_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y127_SLICE_X155Y127_CO5),
.O6(CLBLM_L_X98Y127_SLICE_X155Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y127_SLICE_X155Y127_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y128_SLICE_X154Y128_CQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y127_SLICE_X155Y127_BO5),
.O6(CLBLM_L_X98Y127_SLICE_X155Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0aaa0000aa)
  ) CLBLM_L_X98Y127_SLICE_X155Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y127_SLICE_X154Y127_CO6),
.I3(CLBLM_L_X98Y127_SLICE_X154Y127_B5Q),
.I4(CLBLL_L_X100Y127_SLICE_X157Y127_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y127_SLICE_X155Y127_AO5),
.O6(CLBLM_L_X98Y127_SLICE_X155Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y128_SLICE_X154Y128_AO5),
.Q(CLBLM_L_X98Y128_SLICE_X154Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y128_SLICE_X154Y128_BO5),
.Q(CLBLM_L_X98Y128_SLICE_X154Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y128_SLICE_X154Y128_CO5),
.Q(CLBLM_L_X98Y128_SLICE_X154Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y128_SLICE_X154Y128_AO6),
.Q(CLBLM_L_X98Y128_SLICE_X154Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y128_SLICE_X154Y128_BO6),
.Q(CLBLM_L_X98Y128_SLICE_X154Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y128_SLICE_X154Y128_CO6),
.Q(CLBLM_L_X98Y128_SLICE_X154Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_DLUT (
.I0(CLBLM_L_X98Y128_SLICE_X154Y128_C5Q),
.I1(1'b1),
.I2(CLBLM_L_X98Y128_SLICE_X154Y128_BQ),
.I3(CLBLL_L_X100Y129_SLICE_X157Y129_AQ),
.I4(CLBLM_L_X98Y128_SLICE_X154Y128_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_L_X98Y128_SLICE_X154Y128_DO5),
.O6(CLBLM_L_X98Y128_SLICE_X154Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff000000)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_CLUT (
.I0(CLBLM_R_X101Y128_SLICE_X158Y128_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y128_SLICE_X154Y128_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X154Y128_CO5),
.O6(CLBLM_L_X98Y128_SLICE_X154Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y128_SLICE_X154Y128_BQ),
.I2(CLBLL_L_X100Y129_SLICE_X157Y129_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X154Y128_BO5),
.O6(CLBLM_L_X98Y128_SLICE_X154Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa88882222)
  ) CLBLM_L_X98Y128_SLICE_X154Y128_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y128_SLICE_X154Y128_C5Q),
.I2(1'b1),
.I3(CLBLM_R_X97Y124_SLICE_X152Y124_CO6),
.I4(CLBLM_R_X97Y127_SLICE_X153Y127_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X154Y128_AO5),
.O6(CLBLM_L_X98Y128_SLICE_X154Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y128_SLICE_X155Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X155Y128_DO5),
.O6(CLBLM_L_X98Y128_SLICE_X155Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y128_SLICE_X155Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X155Y128_CO5),
.O6(CLBLM_L_X98Y128_SLICE_X155Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y128_SLICE_X155Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X155Y128_BO5),
.O6(CLBLM_L_X98Y128_SLICE_X155Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y128_SLICE_X155Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y128_SLICE_X155Y128_AO5),
.O6(CLBLM_L_X98Y128_SLICE_X155Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X154Y129_BO5),
.Q(CLBLM_L_X98Y129_SLICE_X154Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X155Y129_BO5),
.Q(CLBLM_L_X98Y129_SLICE_X154Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X154Y129_BO6),
.Q(CLBLM_L_X98Y129_SLICE_X154Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X154Y129_AO5),
.Q(CLBLM_L_X98Y129_SLICE_X154Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y129_SLICE_X154Y129_DO5),
.O6(CLBLM_L_X98Y129_SLICE_X154Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_CLUT (
.I0(CLBLM_L_X98Y129_SLICE_X154Y129_BQ),
.I1(CLBLM_L_X98Y129_SLICE_X154Y129_CQ),
.I2(CLBLM_R_X97Y129_SLICE_X152Y129_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X98Y129_SLICE_X154Y129_B5Q),
.I5(CLBLM_L_X98Y130_SLICE_X155Y130_CQ),
.O5(CLBLM_L_X98Y129_SLICE_X154Y129_CO5),
.O6(CLBLM_L_X98Y129_SLICE_X154Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y129_SLICE_X154Y129_BQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y130_SLICE_X155Y130_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y129_SLICE_X154Y129_BO5),
.O6(CLBLM_L_X98Y129_SLICE_X154Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55a88888888)
  ) CLBLM_L_X98Y129_SLICE_X154Y129_ALUT (
.I0(CLBLM_L_X98Y129_SLICE_X154Y129_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X98Y129_SLICE_X154Y129_CQ),
.I3(CLBLM_L_X98Y130_SLICE_X155Y130_CQ),
.I4(CLBLM_L_X98Y129_SLICE_X154Y129_BQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y129_SLICE_X154Y129_AO5),
.O6(CLBLM_L_X98Y129_SLICE_X154Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X155Y129_AO5),
.Q(CLBLM_L_X98Y129_SLICE_X155Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X155Y129_CO5),
.Q(CLBLM_L_X98Y129_SLICE_X155Y129_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X155Y129_AO6),
.Q(CLBLM_L_X98Y129_SLICE_X155Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y129_SLICE_X155Y129_CO6),
.Q(CLBLM_L_X98Y129_SLICE_X155Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12ed21ed21de12)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_DLUT (
.I0(CLBLM_L_X98Y129_SLICE_X155Y129_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X98Y130_SLICE_X155Y130_BQ),
.I3(CLBLM_R_X97Y130_SLICE_X153Y130_AQ),
.I4(CLBLM_L_X98Y129_SLICE_X154Y129_AQ),
.I5(CLBLM_L_X98Y129_SLICE_X155Y129_CQ),
.O5(CLBLM_L_X98Y129_SLICE_X155Y129_DO5),
.O6(CLBLM_L_X98Y129_SLICE_X155Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_L_X98Y130_SLICE_X155Y130_BQ),
.I4(CLBLM_L_X98Y129_SLICE_X155Y129_CQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y129_SLICE_X155Y129_CO5),
.O6(CLBLM_L_X98Y129_SLICE_X155Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_BLUT (
.I0(CLBLM_L_X98Y129_SLICE_X154Y129_AQ),
.I1(CLBLM_L_X98Y130_SLICE_X155Y130_BQ),
.I2(CLBLM_L_X98Y129_SLICE_X155Y129_CQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y129_SLICE_X155Y129_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y129_SLICE_X155Y129_BO5),
.O6(CLBLM_L_X98Y129_SLICE_X155Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000000f000f00)
  ) CLBLM_L_X98Y129_SLICE_X155Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X98Y129_SLICE_X155Y129_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y127_SLICE_X154Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y129_SLICE_X155Y129_AO5),
.O6(CLBLM_L_X98Y129_SLICE_X155Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X154Y130_BO5),
.Q(CLBLM_L_X98Y130_SLICE_X154Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X154Y130_CO5),
.Q(CLBLM_L_X98Y130_SLICE_X154Y130_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X154Y130_AO6),
.Q(CLBLM_L_X98Y130_SLICE_X154Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X154Y130_CO6),
.Q(CLBLM_L_X98Y130_SLICE_X154Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_DLUT (
.I0(CLBLM_L_X98Y130_SLICE_X154Y130_C5Q),
.I1(CLBLM_L_X98Y130_SLICE_X154Y130_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y130_SLICE_X154Y130_A5Q),
.I4(CLBLM_L_X98Y130_SLICE_X154Y130_CQ),
.I5(CLBLM_R_X97Y129_SLICE_X152Y129_CQ),
.O5(CLBLM_L_X98Y130_SLICE_X154Y130_DO5),
.O6(CLBLM_L_X98Y130_SLICE_X154Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y130_SLICE_X154Y130_CQ),
.I2(CLBLM_L_X98Y130_SLICE_X154Y130_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y130_SLICE_X154Y130_CO5),
.O6(CLBLM_L_X98Y130_SLICE_X154Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y130_SLICE_X154Y130_A5Q),
.I2(CLBLM_L_X98Y130_SLICE_X154Y130_AQ),
.I3(CLBLM_L_X98Y130_SLICE_X154Y130_CQ),
.I4(CLBLM_L_X98Y130_SLICE_X154Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y130_SLICE_X154Y130_BO5),
.O6(CLBLM_L_X98Y130_SLICE_X154Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ee2200000000)
  ) CLBLM_L_X98Y130_SLICE_X154Y130_ALUT (
.I0(CLBLL_L_X102Y130_SLICE_X160Y130_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y133_SLICE_X154Y133_AQ),
.I3(CLBLM_L_X98Y130_SLICE_X154Y130_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y130_SLICE_X154Y130_AO5),
.O6(CLBLM_L_X98Y130_SLICE_X154Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X155Y130_AO5),
.Q(CLBLM_L_X98Y130_SLICE_X155Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X155Y130_DO5),
.Q(CLBLM_L_X98Y130_SLICE_X155Y130_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X155Y130_AO6),
.Q(CLBLM_L_X98Y130_SLICE_X155Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X155Y130_BO6),
.Q(CLBLM_L_X98Y130_SLICE_X155Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X155Y130_CO6),
.Q(CLBLM_L_X98Y130_SLICE_X155Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y130_SLICE_X155Y130_DO6),
.Q(CLBLM_L_X98Y130_SLICE_X155Y130_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8844884448488484)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_DLUT (
.I0(CLBLM_L_X98Y128_SLICE_X154Y128_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X98Y132_SLICE_X155Y132_CQ),
.I3(CLBLM_L_X98Y129_SLICE_X154Y129_CQ),
.I4(CLBLM_R_X97Y130_SLICE_X152Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y130_SLICE_X155Y130_DO5),
.O6(CLBLM_L_X98Y130_SLICE_X155Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8cc000808cc00)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_CLUT (
.I0(CLBLM_L_X98Y129_SLICE_X154Y129_AO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X102Y131_SLICE_X160Y131_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X98Y129_SLICE_X155Y129_A5Q),
.O5(CLBLM_L_X98Y130_SLICE_X155Y130_CO5),
.O6(CLBLM_L_X98Y130_SLICE_X155Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heee22e2200000000)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_BLUT (
.I0(CLBLM_R_X101Y130_SLICE_X159Y130_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y129_SLICE_X155Y129_BO6),
.I4(CLBLM_L_X98Y130_SLICE_X155Y130_A5Q),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y130_SLICE_X155Y130_BO5),
.O6(CLBLM_L_X98Y130_SLICE_X155Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_L_X98Y130_SLICE_X155Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y130_SLICE_X155Y130_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y129_SLICE_X155Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y130_SLICE_X155Y130_AO5),
.O6(CLBLM_L_X98Y130_SLICE_X155Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X154Y131_BO5),
.Q(CLBLM_L_X98Y131_SLICE_X154Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X154Y131_CO5),
.Q(CLBLM_L_X98Y131_SLICE_X154Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.Q(CLBLM_L_X98Y131_SLICE_X154Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X154Y131_CO6),
.Q(CLBLM_L_X98Y131_SLICE_X154Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_DLUT (
.I0(CLBLM_L_X98Y131_SLICE_X154Y131_C5Q),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_CQ),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AQ),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X97Y130_SLICE_X153Y130_A5Q),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_DO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000cccc0000)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_CQ),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_CO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_A5Q),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AQ),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_CQ),
.I4(CLBLM_L_X98Y131_SLICE_X154Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_BO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a82020a820a820)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X101Y131_SLICE_X158Y131_DO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_BO6),
.I4(CLBLM_L_X98Y130_SLICE_X155Y130_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_AO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X155Y131_AO5),
.Q(CLBLM_L_X98Y131_SLICE_X155Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X155Y131_CO5),
.Q(CLBLM_L_X98Y131_SLICE_X155Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X155Y131_DO5),
.Q(CLBLM_L_X98Y131_SLICE_X155Y131_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X155Y131_AO6),
.Q(CLBLM_L_X98Y131_SLICE_X155Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X155Y131_BO6),
.Q(CLBLM_L_X98Y131_SLICE_X155Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y131_SLICE_X155Y131_DO6),
.Q(CLBLM_L_X98Y131_SLICE_X155Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0000aa82828282)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_A5Q),
.I2(CLBLM_L_X98Y131_SLICE_X155Y131_DQ),
.I3(CLBLM_L_X98Y129_SLICE_X154Y129_AQ),
.I4(CLBLM_L_X98Y130_SLICE_X155Y130_DQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_DO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966c0c0c0c0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_CLUT (
.I0(CLBLM_R_X97Y131_SLICE_X153Y131_BQ),
.I1(CLBLM_R_X97Y131_SLICE_X153Y131_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y132_SLICE_X155Y132_BQ),
.I4(CLBLM_L_X98Y131_SLICE_X155Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_CO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0bb8800000000)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_BLUT (
.I0(CLBLM_R_X97Y130_SLICE_X152Y130_AO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y131_SLICE_X155Y131_AQ),
.I3(CLBLM_R_X101Y132_SLICE_X159Y132_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_BO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y131_SLICE_X155Y131_A5Q),
.I2(CLBLM_L_X98Y130_SLICE_X155Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_AO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X154Y132_BO5),
.Q(CLBLM_L_X98Y132_SLICE_X154Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X154Y132_CO5),
.Q(CLBLM_L_X98Y132_SLICE_X154Y132_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.Q(CLBLM_L_X98Y132_SLICE_X154Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X154Y132_CO6),
.Q(CLBLM_L_X98Y132_SLICE_X154Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_DLUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X98Y132_SLICE_X154Y132_AQ),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_A5Q),
.I4(CLBLM_R_X97Y132_SLICE_X153Y132_CQ),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_CQ),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_DO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X98Y132_SLICE_X154Y132_CQ),
.I2(CLBLM_L_X98Y132_SLICE_X154Y132_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_CO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y132_SLICE_X154Y132_A5Q),
.I2(CLBLM_L_X98Y132_SLICE_X154Y132_AQ),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_CQ),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_BO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88f0f000000000)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X98Y133_SLICE_X154Y133_BQ),
.I2(CLBLM_R_X101Y133_SLICE_X159Y133_BO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_AO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X155Y132_CO5),
.Q(CLBLM_L_X98Y132_SLICE_X155Y132_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X155Y132_AO5),
.Q(CLBLM_L_X98Y132_SLICE_X155Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X155Y132_BO6),
.Q(CLBLM_L_X98Y132_SLICE_X155Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y132_SLICE_X155Y132_CO6),
.Q(CLBLM_L_X98Y132_SLICE_X155Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_DO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00cc00c88884444)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_CLUT (
.I0(CLBLM_L_X98Y130_SLICE_X155Y130_D5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X98Y131_SLICE_X155Y131_B5Q),
.I3(CLBLM_L_X98Y131_SLICE_X155Y131_D5Q),
.I4(CLBLM_L_X98Y132_SLICE_X155Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_CO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbc83b0800000000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_BLUT (
.I0(CLBLM_L_X98Y131_SLICE_X155Y131_CO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X101Y133_SLICE_X158Y133_DO6),
.I4(CLBLM_L_X98Y131_SLICE_X155Y131_A5Q),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_BO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f000f000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_ALUT (
.I0(CLBLM_L_X98Y133_SLICE_X155Y133_BQ),
.I1(CLBLM_R_X97Y132_SLICE_X153Y132_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y132_SLICE_X153Y132_A5Q),
.I4(CLBLM_L_X98Y132_SLICE_X155Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_AO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X154Y133_AO5),
.Q(CLBLM_L_X98Y133_SLICE_X154Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X154Y133_BO5),
.Q(CLBLM_L_X98Y133_SLICE_X154Y133_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X154Y133_AO6),
.Q(CLBLM_L_X98Y133_SLICE_X154Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X154Y133_BO6),
.Q(CLBLM_L_X98Y133_SLICE_X154Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X154Y133_DO5),
.O6(CLBLM_L_X98Y133_SLICE_X154Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X154Y133_CO5),
.O6(CLBLM_L_X98Y133_SLICE_X154Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaaa0000)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y133_SLICE_X154Y133_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y133_SLICE_X155Y133_AQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X154Y133_BO5),
.O6(CLBLM_L_X98Y133_SLICE_X154Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X98Y133_SLICE_X154Y133_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y133_SLICE_X154Y133_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y133_SLICE_X154Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X154Y133_AO5),
.O6(CLBLM_L_X98Y133_SLICE_X154Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X155Y133_AO5),
.Q(CLBLM_L_X98Y133_SLICE_X155Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X155Y133_AO6),
.Q(CLBLM_L_X98Y133_SLICE_X155Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y133_SLICE_X155Y133_BO6),
.Q(CLBLM_L_X98Y133_SLICE_X155Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X155Y133_DO5),
.O6(CLBLM_L_X98Y133_SLICE_X155Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X155Y133_CO5),
.O6(CLBLM_L_X98Y133_SLICE_X155Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8ad58000000000)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X98Y133_SLICE_X155Y133_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y134_SLICE_X156Y134_CO6),
.I4(CLBLM_L_X98Y132_SLICE_X155Y132_AO6),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y133_SLICE_X155Y133_BO5),
.O6(CLBLM_L_X98Y133_SLICE_X155Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_L_X98Y133_SLICE_X155Y133_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y133_SLICE_X155Y133_A5Q),
.I2(CLBLM_L_X98Y131_SLICE_X155Y131_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y133_SLICE_X155Y133_AO5),
.O6(CLBLM_L_X98Y133_SLICE_X155Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y134_SLICE_X154Y134_BO5),
.Q(CLBLM_L_X98Y134_SLICE_X154Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y134_SLICE_X154Y134_CO5),
.Q(CLBLM_L_X98Y134_SLICE_X154Y134_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y134_SLICE_X154Y134_AO6),
.Q(CLBLM_L_X98Y134_SLICE_X154Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_L_X98Y134_SLICE_X154Y134_CO6),
.Q(CLBLM_L_X98Y134_SLICE_X154Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_DLUT (
.I0(CLBLM_L_X98Y134_SLICE_X154Y134_C5Q),
.I1(CLBLM_L_X98Y134_SLICE_X154Y134_AQ),
.I2(CLBLM_R_X97Y132_SLICE_X153Y132_B5Q),
.I3(CLBLM_L_X98Y134_SLICE_X154Y134_A5Q),
.I4(CLBLM_L_X98Y134_SLICE_X154Y134_CQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_L_X98Y134_SLICE_X154Y134_DO5),
.O6(CLBLM_L_X98Y134_SLICE_X154Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff000000)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X98Y134_SLICE_X154Y134_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y134_SLICE_X154Y134_CQ),
.I5(1'b1),
.O5(CLBLM_L_X98Y134_SLICE_X154Y134_CO5),
.O6(CLBLM_L_X98Y134_SLICE_X154Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_BLUT (
.I0(CLBLM_L_X98Y134_SLICE_X154Y134_CQ),
.I1(CLBLM_L_X98Y134_SLICE_X154Y134_A5Q),
.I2(CLBLM_L_X98Y134_SLICE_X154Y134_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X98Y134_SLICE_X154Y134_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X98Y134_SLICE_X154Y134_BO5),
.O6(CLBLM_L_X98Y134_SLICE_X154Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cccc00000000)
  ) CLBLM_L_X98Y134_SLICE_X154Y134_ALUT (
.I0(CLBLM_L_X98Y133_SLICE_X154Y133_B5Q),
.I1(CLBLL_L_X102Y135_SLICE_X160Y135_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y134_SLICE_X154Y134_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_L_X98Y134_SLICE_X154Y134_AO5),
.O6(CLBLM_L_X98Y134_SLICE_X154Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y134_SLICE_X155Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y134_SLICE_X155Y134_DO5),
.O6(CLBLM_L_X98Y134_SLICE_X155Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y134_SLICE_X155Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y134_SLICE_X155Y134_CO5),
.O6(CLBLM_L_X98Y134_SLICE_X155Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y134_SLICE_X155Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y134_SLICE_X155Y134_BO5),
.O6(CLBLM_L_X98Y134_SLICE_X155Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y134_SLICE_X155Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y134_SLICE_X155Y134_AO5),
.O6(CLBLM_L_X98Y134_SLICE_X155Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y114_SLICE_X140Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X140Y114_DO5),
.O6(CLBLM_R_X89Y114_SLICE_X140Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y114_SLICE_X140Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X140Y114_CO5),
.O6(CLBLM_R_X89Y114_SLICE_X140Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y114_SLICE_X140Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X140Y114_BO5),
.O6(CLBLM_R_X89Y114_SLICE_X140Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y114_SLICE_X140Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X140Y114_AO5),
.O6(CLBLM_R_X89Y114_SLICE_X140Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y114_SLICE_X141Y114_AO5),
.Q(CLBLM_R_X89Y114_SLICE_X141Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y114_SLICE_X141Y114_BO5),
.Q(CLBLM_R_X89Y114_SLICE_X141Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y114_SLICE_X141Y114_AO6),
.Q(CLBLM_R_X89Y114_SLICE_X141Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y114_SLICE_X141Y114_BO6),
.Q(CLBLM_R_X89Y114_SLICE_X141Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X141Y114_DO5),
.O6(CLBLM_R_X89Y114_SLICE_X141Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X89Y114_SLICE_X141Y114_BQ),
.I3(CLBLM_L_X90Y116_SLICE_X143Y116_BQ),
.I4(CLBLM_R_X89Y114_SLICE_X141Y114_B5Q),
.I5(CLBLM_R_X89Y114_SLICE_X141Y114_AQ),
.O5(CLBLM_R_X89Y114_SLICE_X141Y114_CO5),
.O6(CLBLM_R_X89Y114_SLICE_X141Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y114_SLICE_X141Y114_AQ),
.I3(1'b1),
.I4(CLBLM_R_X89Y114_SLICE_X141Y114_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X141Y114_BO5),
.O6(CLBLM_R_X89Y114_SLICE_X141Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X89Y114_SLICE_X141Y114_ALUT (
.I0(CLBLM_L_X90Y116_SLICE_X143Y116_BQ),
.I1(CLBLM_L_X90Y114_SLICE_X142Y114_C5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y114_SLICE_X141Y114_AO5),
.O6(CLBLM_R_X89Y114_SLICE_X141Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X140Y115_BO5),
.Q(CLBLM_R_X89Y115_SLICE_X140Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X140Y115_CO5),
.Q(CLBLM_R_X89Y115_SLICE_X140Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X140Y115_AO6),
.Q(CLBLM_R_X89Y115_SLICE_X140Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X140Y115_CO6),
.Q(CLBLM_R_X89Y115_SLICE_X140Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_DLUT (
.I0(CLBLM_R_X89Y115_SLICE_X140Y115_C5Q),
.I1(CLBLM_R_X89Y115_SLICE_X140Y115_CQ),
.I2(CLBLM_R_X89Y115_SLICE_X140Y115_AQ),
.I3(CLBLM_R_X89Y115_SLICE_X140Y115_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y116_SLICE_X141Y116_C5Q),
.O5(CLBLM_R_X89Y115_SLICE_X140Y115_DO5),
.O6(CLBLM_R_X89Y115_SLICE_X140Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y115_SLICE_X140Y115_CQ),
.I2(CLBLM_R_X89Y115_SLICE_X140Y115_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y115_SLICE_X140Y115_CO5),
.O6(CLBLM_R_X89Y115_SLICE_X140Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_BLUT (
.I0(CLBLM_R_X89Y115_SLICE_X140Y115_CQ),
.I1(CLBLM_R_X89Y115_SLICE_X140Y115_A5Q),
.I2(CLBLM_R_X89Y115_SLICE_X140Y115_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X89Y115_SLICE_X140Y115_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y115_SLICE_X140Y115_BO5),
.O6(CLBLM_R_X89Y115_SLICE_X140Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cccc00000000)
  ) CLBLM_R_X89Y115_SLICE_X140Y115_ALUT (
.I0(CLBLM_R_X89Y116_SLICE_X140Y116_A5Q),
.I1(CLBLM_L_X90Y119_SLICE_X143Y119_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X89Y115_SLICE_X140Y115_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X89Y115_SLICE_X140Y115_AO5),
.O6(CLBLM_R_X89Y115_SLICE_X140Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X141Y115_AO5),
.Q(CLBLM_R_X89Y115_SLICE_X141Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X141Y115_BO5),
.Q(CLBLM_R_X89Y115_SLICE_X141Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X141Y115_AO6),
.Q(CLBLM_R_X89Y115_SLICE_X141Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X141Y115_BO6),
.Q(CLBLM_R_X89Y115_SLICE_X141Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y115_SLICE_X141Y115_CO6),
.Q(CLBLM_R_X89Y115_SLICE_X141Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_DLUT (
.I0(CLBLM_L_X90Y115_SLICE_X142Y115_AQ),
.I1(CLBLM_R_X89Y115_SLICE_X141Y115_AQ),
.I2(1'b1),
.I3(CLBLM_R_X89Y115_SLICE_X141Y115_A5Q),
.I4(CLBLM_R_X89Y115_SLICE_X141Y115_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X89Y115_SLICE_X141Y115_DO5),
.O6(CLBLM_R_X89Y115_SLICE_X141Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4488884444888844)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_CLUT (
.I0(CLBLM_R_X89Y116_SLICE_X141Y116_C5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y117_SLICE_X146Y117_A5Q),
.I4(CLBLM_R_X89Y115_SLICE_X141Y115_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y115_SLICE_X141Y115_CO5),
.O6(CLBLM_R_X89Y115_SLICE_X141Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00c0c0c0c0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y115_SLICE_X141Y115_A5Q),
.I3(CLBLM_R_X89Y118_SLICE_X141Y118_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y115_SLICE_X141Y115_BO5),
.O6(CLBLM_R_X89Y115_SLICE_X141Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00c0c0c0c0)
  ) CLBLM_R_X89Y115_SLICE_X141Y115_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y115_SLICE_X141Y115_AQ),
.I3(CLBLM_L_X90Y115_SLICE_X142Y115_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y115_SLICE_X141Y115_AO5),
.O6(CLBLM_R_X89Y115_SLICE_X141Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X140Y116_AO5),
.Q(CLBLM_R_X89Y116_SLICE_X140Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X141Y116_AO5),
.Q(CLBLM_R_X89Y116_SLICE_X140Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X140Y116_AO6),
.Q(CLBLM_R_X89Y116_SLICE_X140Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X140Y116_BO6),
.Q(CLBLM_R_X89Y116_SLICE_X140Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y116_SLICE_X140Y116_DO5),
.O6(CLBLM_R_X89Y116_SLICE_X140Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y116_SLICE_X140Y116_CO5),
.O6(CLBLM_R_X89Y116_SLICE_X140Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8ccc80040cc4000)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y116_SLICE_X141Y116_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X90Y120_SLICE_X142Y120_DO6),
.I5(CLBLM_R_X89Y117_SLICE_X140Y117_CQ),
.O5(CLBLM_R_X89Y116_SLICE_X140Y116_BO5),
.O6(CLBLM_R_X89Y116_SLICE_X140Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X89Y116_SLICE_X140Y116_ALUT (
.I0(CLBLM_R_X89Y117_SLICE_X140Y117_CQ),
.I1(CLBLM_R_X89Y116_SLICE_X140Y116_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y116_SLICE_X140Y116_AO5),
.O6(CLBLM_R_X89Y116_SLICE_X140Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X141Y116_BO5),
.Q(CLBLM_R_X89Y116_SLICE_X141Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X141Y116_CO5),
.Q(CLBLM_R_X89Y116_SLICE_X141Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X141Y116_BO6),
.Q(CLBLM_R_X89Y116_SLICE_X141Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y116_SLICE_X141Y116_CO6),
.Q(CLBLM_R_X89Y116_SLICE_X141Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc5acca5cca5cc5a)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_DLUT (
.I0(CLBLM_R_X89Y116_SLICE_X141Y116_BQ),
.I1(CLBLM_R_X89Y116_SLICE_X141Y116_CQ),
.I2(CLBLM_R_X89Y116_SLICE_X140Y116_B5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X89Y116_SLICE_X141Y116_B5Q),
.I5(CLBLM_R_X89Y116_SLICE_X140Y116_BQ),
.O5(CLBLM_R_X89Y116_SLICE_X141Y116_DO5),
.O6(CLBLM_R_X89Y116_SLICE_X141Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_CLUT (
.I0(CLBLM_L_X90Y116_SLICE_X142Y116_BQ),
.I1(CLBLM_R_X89Y116_SLICE_X141Y116_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y117_SLICE_X142Y117_A5Q),
.I4(CLBLM_R_X89Y118_SLICE_X141Y118_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y116_SLICE_X141Y116_CO5),
.O6(CLBLM_R_X89Y116_SLICE_X141Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X89Y116_SLICE_X140Y116_BQ),
.I4(CLBLM_R_X89Y116_SLICE_X141Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y116_SLICE_X141Y116_BO5),
.O6(CLBLM_R_X89Y116_SLICE_X141Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_R_X89Y116_SLICE_X141Y116_ALUT (
.I0(CLBLM_R_X89Y116_SLICE_X141Y116_B5Q),
.I1(CLBLM_R_X89Y116_SLICE_X141Y116_BQ),
.I2(CLBLM_R_X89Y116_SLICE_X140Y116_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X89Y116_SLICE_X140Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y116_SLICE_X141Y116_AO5),
.O6(CLBLM_R_X89Y116_SLICE_X141Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X140Y117_AO5),
.Q(CLBLM_R_X89Y117_SLICE_X140Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X140Y117_CO5),
.Q(CLBLM_R_X89Y117_SLICE_X140Y117_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X140Y117_AO6),
.Q(CLBLM_R_X89Y117_SLICE_X140Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X140Y117_BO6),
.Q(CLBLM_R_X89Y117_SLICE_X140Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X140Y117_CO6),
.Q(CLBLM_R_X89Y117_SLICE_X140Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y117_SLICE_X140Y117_DO5),
.O6(CLBLM_R_X89Y117_SLICE_X140Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y119_SLICE_X140Y119_BQ),
.I2(CLBLM_R_X89Y117_SLICE_X140Y117_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y117_SLICE_X140Y117_CO5),
.O6(CLBLM_R_X89Y117_SLICE_X140Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc000c088c088c0)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_BLUT (
.I0(CLBLM_L_X90Y119_SLICE_X142Y119_AO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y117_SLICE_X141Y117_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X89Y118_SLICE_X140Y118_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y117_SLICE_X140Y117_BO5),
.O6(CLBLM_R_X89Y117_SLICE_X140Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X89Y117_SLICE_X140Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y117_SLICE_X140Y117_A5Q),
.I2(CLBLM_R_X89Y118_SLICE_X140Y118_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y117_SLICE_X140Y117_AO5),
.O6(CLBLM_R_X89Y117_SLICE_X140Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X141Y117_BO5),
.Q(CLBLM_R_X89Y117_SLICE_X141Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X141Y117_CO5),
.Q(CLBLM_R_X89Y117_SLICE_X141Y117_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X141Y117_AO6),
.Q(CLBLM_R_X89Y117_SLICE_X141Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y117_SLICE_X141Y117_CO6),
.Q(CLBLM_R_X89Y117_SLICE_X141Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0069699696)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_DLUT (
.I0(CLBLM_R_X89Y117_SLICE_X141Y117_C5Q),
.I1(CLBLM_R_X89Y117_SLICE_X141Y117_CQ),
.I2(CLBLM_R_X89Y117_SLICE_X141Y117_A5Q),
.I3(CLBLM_R_X89Y118_SLICE_X141Y118_D5Q),
.I4(CLBLM_R_X89Y117_SLICE_X141Y117_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y117_SLICE_X141Y117_DO5),
.O6(CLBLM_R_X89Y117_SLICE_X141Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y117_SLICE_X141Y117_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X89Y117_SLICE_X141Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y117_SLICE_X141Y117_CO5),
.O6(CLBLM_R_X89Y117_SLICE_X141Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_BLUT (
.I0(CLBLM_R_X89Y117_SLICE_X141Y117_CQ),
.I1(CLBLM_R_X89Y117_SLICE_X141Y117_A5Q),
.I2(CLBLM_R_X89Y117_SLICE_X141Y117_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X89Y117_SLICE_X141Y117_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y117_SLICE_X141Y117_BO5),
.O6(CLBLM_R_X89Y117_SLICE_X141Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he200e200ee002200)
  ) CLBLM_R_X89Y117_SLICE_X141Y117_ALUT (
.I0(CLBLM_R_X89Y120_SLICE_X141Y120_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X89Y117_SLICE_X140Y117_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X89Y117_SLICE_X141Y117_BO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y117_SLICE_X141Y117_AO5),
.O6(CLBLM_R_X89Y117_SLICE_X141Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X140Y118_AO5),
.Q(CLBLM_R_X89Y118_SLICE_X140Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X140Y118_CO5),
.Q(CLBLM_R_X89Y118_SLICE_X140Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X140Y118_DO5),
.Q(CLBLM_R_X89Y118_SLICE_X140Y118_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X140Y118_AO6),
.Q(CLBLM_R_X89Y118_SLICE_X140Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X140Y118_BO6),
.Q(CLBLM_R_X89Y118_SLICE_X140Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X140Y118_DO6),
.Q(CLBLM_R_X89Y118_SLICE_X140Y118_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X92Y122_SLICE_X145Y122_BQ),
.I3(1'b1),
.I4(CLBLM_R_X89Y118_SLICE_X140Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y118_SLICE_X140Y118_DO5),
.O6(CLBLM_R_X89Y118_SLICE_X140Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caa00aa00)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y118_SLICE_X140Y118_B5Q),
.I2(CLBLM_R_X89Y118_SLICE_X140Y118_DQ),
.I3(CLBLM_L_X90Y118_SLICE_X142Y118_A5Q),
.I4(CLBLM_R_X89Y118_SLICE_X140Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y118_SLICE_X140Y118_CO5),
.O6(CLBLM_R_X89Y118_SLICE_X140Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd000008f800000)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X89Y118_SLICE_X140Y118_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_R_X87Y118_SLICE_X139Y118_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X89Y118_SLICE_X140Y118_CO6),
.O5(CLBLM_R_X89Y118_SLICE_X140Y118_BO5),
.O6(CLBLM_R_X89Y118_SLICE_X140Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f0f00000)
  ) CLBLM_R_X89Y118_SLICE_X140Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y118_SLICE_X140Y118_A5Q),
.I2(CLBLM_R_X89Y119_SLICE_X140Y119_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X89Y118_SLICE_X140Y118_AO5),
.O6(CLBLM_R_X89Y118_SLICE_X140Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X141Y118_BO5),
.Q(CLBLM_R_X89Y118_SLICE_X141Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X141Y118_DO5),
.Q(CLBLM_R_X89Y118_SLICE_X141Y118_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X141Y118_AO6),
.Q(CLBLM_R_X89Y118_SLICE_X141Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X141Y118_CO6),
.Q(CLBLM_R_X89Y118_SLICE_X141Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y118_SLICE_X141Y118_DO6),
.Q(CLBLM_R_X89Y118_SLICE_X141Y118_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc330000a5a50000)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_DLUT (
.I0(CLBLM_L_X90Y119_SLICE_X143Y119_AQ),
.I1(CLBLM_R_X89Y118_SLICE_X141Y118_CQ),
.I2(CLBLM_R_X89Y118_SLICE_X141Y118_DQ),
.I3(CLBLM_R_X89Y118_SLICE_X140Y118_B5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X89Y118_SLICE_X141Y118_DO5),
.O6(CLBLM_R_X89Y118_SLICE_X141Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2288882222888822)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y117_SLICE_X146Y117_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X89Y118_SLICE_X141Y118_A5Q),
.I4(CLBLM_R_X89Y120_SLICE_X140Y120_CQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y118_SLICE_X141Y118_CO5),
.O6(CLBLM_R_X89Y118_SLICE_X141Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_BLUT (
.I0(CLBLM_L_X92Y118_SLICE_X144Y118_A5Q),
.I1(CLBLM_R_X89Y118_SLICE_X141Y118_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y115_SLICE_X141Y115_BQ),
.I4(CLBLM_R_X89Y118_SLICE_X141Y118_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y118_SLICE_X141Y118_BO5),
.O6(CLBLM_R_X89Y118_SLICE_X141Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e02020e020e020)
  ) CLBLM_R_X89Y118_SLICE_X141Y118_ALUT (
.I0(CLBLM_R_X89Y119_SLICE_X141Y119_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y118_SLICE_X141Y118_BO6),
.I4(CLBLM_R_X89Y119_SLICE_X140Y119_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y118_SLICE_X141Y118_AO5),
.O6(CLBLM_R_X89Y118_SLICE_X141Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X140Y119_AO5),
.Q(CLBLM_R_X89Y119_SLICE_X140Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X140Y119_BO5),
.Q(CLBLM_R_X89Y119_SLICE_X140Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X140Y119_AO6),
.Q(CLBLM_R_X89Y119_SLICE_X140Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X140Y119_BO6),
.Q(CLBLM_R_X89Y119_SLICE_X140Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y119_SLICE_X140Y119_DO5),
.O6(CLBLM_R_X89Y119_SLICE_X140Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y119_SLICE_X140Y119_CO5),
.O6(CLBLM_R_X89Y119_SLICE_X140Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0c0c0c0)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_BLUT (
.I0(CLBLM_R_X89Y119_SLICE_X140Y119_B5Q),
.I1(CLBLM_R_X89Y124_SLICE_X140Y124_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y119_SLICE_X140Y119_BO5),
.O6(CLBLM_R_X89Y119_SLICE_X140Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_R_X89Y119_SLICE_X140Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y119_SLICE_X140Y119_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X92Y123_SLICE_X145Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y119_SLICE_X140Y119_AO5),
.O6(CLBLM_R_X89Y119_SLICE_X140Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X141Y119_BO5),
.Q(CLBLM_R_X89Y119_SLICE_X141Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X141Y119_CO5),
.Q(CLBLM_R_X89Y119_SLICE_X141Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X141Y119_AO6),
.Q(CLBLM_R_X89Y119_SLICE_X141Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y119_SLICE_X141Y119_CO6),
.Q(CLBLM_R_X89Y119_SLICE_X141Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_DLUT (
.I0(CLBLM_R_X89Y119_SLICE_X141Y119_C5Q),
.I1(CLBLM_R_X89Y119_SLICE_X141Y119_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X89Y119_SLICE_X141Y119_A5Q),
.I4(CLBLM_R_X89Y119_SLICE_X141Y119_AQ),
.I5(CLBLM_R_X89Y118_SLICE_X141Y118_CQ),
.O5(CLBLM_R_X89Y119_SLICE_X141Y119_DO5),
.O6(CLBLM_R_X89Y119_SLICE_X141Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y119_SLICE_X141Y119_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X89Y119_SLICE_X141Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y119_SLICE_X141Y119_CO5),
.O6(CLBLM_R_X89Y119_SLICE_X141Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_BLUT (
.I0(CLBLM_R_X89Y119_SLICE_X141Y119_AQ),
.I1(CLBLM_R_X89Y119_SLICE_X141Y119_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y119_SLICE_X141Y119_CQ),
.I4(CLBLM_R_X89Y119_SLICE_X141Y119_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y119_SLICE_X141Y119_BO5),
.O6(CLBLM_R_X89Y119_SLICE_X141Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d07050a0802000)
  ) CLBLM_R_X89Y119_SLICE_X141Y119_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y119_SLICE_X141Y119_BO6),
.I4(CLBLM_R_X89Y119_SLICE_X140Y119_B5Q),
.I5(CLBLM_L_X90Y122_SLICE_X143Y122_DO6),
.O5(CLBLM_R_X89Y119_SLICE_X141Y119_AO5),
.O6(CLBLM_R_X89Y119_SLICE_X141Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X140Y120_BO5),
.Q(CLBLM_R_X89Y120_SLICE_X140Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X140Y120_AO6),
.Q(CLBLM_R_X89Y120_SLICE_X140Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X140Y120_CO6),
.Q(CLBLM_R_X89Y120_SLICE_X140Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_DLUT (
.I0(CLBLM_L_X92Y122_SLICE_X145Y122_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X89Y120_SLICE_X140Y120_AQ),
.I3(CLBLM_R_X89Y120_SLICE_X140Y120_A5Q),
.I4(CLBLM_R_X89Y118_SLICE_X140Y118_D5Q),
.I5(CLBLM_R_X97Y120_SLICE_X152Y120_BQ),
.O5(CLBLM_R_X89Y120_SLICE_X140Y120_DO5),
.O6(CLBLM_R_X89Y120_SLICE_X140Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0000aaaa0000aa)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X89Y120_SLICE_X140Y120_A5Q),
.I4(CLBLM_L_X92Y123_SLICE_X144Y123_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y120_SLICE_X140Y120_CO5),
.O6(CLBLM_R_X89Y120_SLICE_X140Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966a0a0a0a0)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_BLUT (
.I0(CLBLM_R_X89Y118_SLICE_X140Y118_D5Q),
.I1(CLBLM_L_X92Y122_SLICE_X145Y122_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y120_SLICE_X140Y120_AQ),
.I4(CLBLM_R_X89Y120_SLICE_X140Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y120_SLICE_X140Y120_BO5),
.O6(CLBLM_R_X89Y120_SLICE_X140Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e02020e020e020)
  ) CLBLM_R_X89Y120_SLICE_X140Y120_ALUT (
.I0(CLBLM_R_X89Y121_SLICE_X140Y121_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y120_SLICE_X140Y120_BO6),
.I4(CLBLM_R_X89Y119_SLICE_X140Y119_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y120_SLICE_X140Y120_AO5),
.O6(CLBLM_R_X89Y120_SLICE_X140Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X141Y120_AO5),
.Q(CLBLM_R_X89Y120_SLICE_X141Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X141Y120_CO5),
.Q(CLBLM_R_X89Y120_SLICE_X141Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X141Y120_AO6),
.Q(CLBLM_R_X89Y120_SLICE_X141Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X141Y120_BO6),
.Q(CLBLM_R_X89Y120_SLICE_X141Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y120_SLICE_X141Y120_CO6),
.Q(CLBLM_R_X89Y120_SLICE_X141Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3cc3aaaac33c)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_DLUT (
.I0(CLBLM_R_X89Y120_SLICE_X141Y120_C5Q),
.I1(CLBLM_R_X89Y121_SLICE_X141Y121_A5Q),
.I2(CLBLM_R_X89Y121_SLICE_X141Y121_CQ),
.I3(CLBLM_R_X89Y120_SLICE_X141Y120_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y121_SLICE_X141Y121_AQ),
.O5(CLBLM_R_X89Y120_SLICE_X141Y120_DO5),
.O6(CLBLM_R_X89Y120_SLICE_X141Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00aa00a88882222)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y120_SLICE_X141Y120_CQ),
.I2(CLBLL_R_X87Y118_SLICE_X138Y118_AQ),
.I3(CLBLM_R_X89Y120_SLICE_X141Y120_BQ),
.I4(CLBLM_R_X89Y117_SLICE_X141Y117_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y120_SLICE_X141Y120_CO5),
.O6(CLBLM_R_X89Y120_SLICE_X141Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6060606090909090)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_BLUT (
.I0(CLBLM_R_X89Y124_SLICE_X140Y124_CQ),
.I1(CLBLM_R_X89Y119_SLICE_X141Y119_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X90Y115_SLICE_X142Y115_A5Q),
.O5(CLBLM_R_X89Y120_SLICE_X141Y120_BO5),
.O6(CLBLM_R_X89Y120_SLICE_X141Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_R_X89Y120_SLICE_X141Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y121_SLICE_X141Y121_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y120_SLICE_X142Y120_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y120_SLICE_X141Y120_AO5),
.O6(CLBLM_R_X89Y120_SLICE_X141Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X140Y121_BO5),
.Q(CLBLM_R_X89Y121_SLICE_X140Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X140Y121_CO5),
.Q(CLBLM_R_X89Y121_SLICE_X140Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X140Y121_AO6),
.Q(CLBLM_R_X89Y121_SLICE_X140Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X140Y121_CO6),
.Q(CLBLM_R_X89Y121_SLICE_X140Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_DLUT (
.I0(CLBLM_R_X89Y121_SLICE_X140Y121_C5Q),
.I1(CLBLM_R_X89Y121_SLICE_X140Y121_CQ),
.I2(CLBLM_R_X89Y121_SLICE_X140Y121_AQ),
.I3(CLBLM_R_X89Y121_SLICE_X140Y121_A5Q),
.I4(CLBLM_R_X89Y120_SLICE_X140Y120_CQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y121_SLICE_X140Y121_DO5),
.O6(CLBLM_R_X89Y121_SLICE_X140Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y121_SLICE_X140Y121_CQ),
.I2(CLBLM_R_X89Y121_SLICE_X140Y121_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y121_SLICE_X140Y121_CO5),
.O6(CLBLM_R_X89Y121_SLICE_X140Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_BLUT (
.I0(CLBLM_R_X89Y121_SLICE_X140Y121_AQ),
.I1(CLBLM_R_X89Y121_SLICE_X140Y121_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y121_SLICE_X140Y121_CQ),
.I4(CLBLM_R_X89Y121_SLICE_X140Y121_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y121_SLICE_X140Y121_BO5),
.O6(CLBLM_R_X89Y121_SLICE_X140Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0a0a0f000a0a0)
  ) CLBLM_R_X89Y121_SLICE_X140Y121_ALUT (
.I0(CLBLM_R_X89Y124_SLICE_X140Y124_DO6),
.I1(CLBLM_R_X89Y124_SLICE_X140Y124_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y121_SLICE_X140Y121_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y121_SLICE_X140Y121_AO5),
.O6(CLBLM_R_X89Y121_SLICE_X140Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X141Y121_BO5),
.Q(CLBLM_R_X89Y121_SLICE_X141Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X141Y121_CO5),
.Q(CLBLM_R_X89Y121_SLICE_X141Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X141Y121_AO6),
.Q(CLBLM_R_X89Y121_SLICE_X141Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y121_SLICE_X141Y121_CO6),
.Q(CLBLM_R_X89Y121_SLICE_X141Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_DLUT (
.I0(CLBLM_R_X89Y121_SLICE_X141Y121_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X89Y122_SLICE_X141Y122_BQ),
.I3(CLBLM_R_X89Y122_SLICE_X141Y122_DQ),
.I4(CLBLM_R_X89Y122_SLICE_X141Y122_B5Q),
.I5(CLBLM_R_X89Y120_SLICE_X141Y120_CQ),
.O5(CLBLM_R_X89Y121_SLICE_X141Y121_DO5),
.O6(CLBLM_R_X89Y121_SLICE_X141Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y122_SLICE_X141Y122_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X89Y121_SLICE_X141Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y121_SLICE_X141Y121_CO5),
.O6(CLBLM_R_X89Y121_SLICE_X141Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f000f000)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_BLUT (
.I0(CLBLM_R_X89Y121_SLICE_X141Y121_AQ),
.I1(CLBLM_R_X89Y121_SLICE_X141Y121_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y120_SLICE_X141Y120_A5Q),
.I4(CLBLM_R_X89Y121_SLICE_X141Y121_CQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y121_SLICE_X141Y121_BO5),
.O6(CLBLM_R_X89Y121_SLICE_X141Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e20000ee220000)
  ) CLBLM_R_X89Y121_SLICE_X141Y121_ALUT (
.I0(CLBLM_R_X93Y125_SLICE_X146Y125_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X89Y122_SLICE_X141Y122_AQ),
.I3(CLBLM_R_X89Y121_SLICE_X141Y121_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y121_SLICE_X141Y121_AO5),
.O6(CLBLM_R_X89Y121_SLICE_X141Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X140Y122_BO5),
.Q(CLBLM_R_X89Y122_SLICE_X140Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X140Y122_CO5),
.Q(CLBLM_R_X89Y122_SLICE_X140Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X140Y122_AO6),
.Q(CLBLM_R_X89Y122_SLICE_X140Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X140Y122_CO6),
.Q(CLBLM_R_X89Y122_SLICE_X140Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_DLUT (
.I0(CLBLM_R_X89Y122_SLICE_X140Y122_C5Q),
.I1(CLBLM_R_X89Y122_SLICE_X140Y122_AQ),
.I2(CLBLM_L_X92Y121_SLICE_X145Y121_C5Q),
.I3(CLBLM_R_X89Y122_SLICE_X140Y122_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y122_SLICE_X140Y122_CQ),
.O5(CLBLM_R_X89Y122_SLICE_X140Y122_DO5),
.O6(CLBLM_R_X89Y122_SLICE_X140Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y122_SLICE_X140Y122_CQ),
.I2(CLBLM_R_X89Y122_SLICE_X140Y122_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y122_SLICE_X140Y122_CO5),
.O6(CLBLM_R_X89Y122_SLICE_X140Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_BLUT (
.I0(CLBLM_R_X89Y122_SLICE_X140Y122_AQ),
.I1(CLBLM_R_X89Y122_SLICE_X140Y122_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y122_SLICE_X140Y122_CQ),
.I4(CLBLM_R_X89Y122_SLICE_X140Y122_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y122_SLICE_X140Y122_BO5),
.O6(CLBLM_R_X89Y122_SLICE_X140Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d0a08070502000)
  ) CLBLM_R_X89Y122_SLICE_X140Y122_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y122_SLICE_X140Y122_BO6),
.I4(CLBLM_R_X89Y126_SLICE_X141Y126_DO6),
.I5(CLBLM_L_X90Y121_SLICE_X142Y121_AQ),
.O5(CLBLM_R_X89Y122_SLICE_X140Y122_AO5),
.O6(CLBLM_R_X89Y122_SLICE_X140Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X141Y122_AO5),
.Q(CLBLM_R_X89Y122_SLICE_X141Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X141Y122_CO5),
.Q(CLBLM_R_X89Y122_SLICE_X141Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X141Y122_DO5),
.Q(CLBLM_R_X89Y122_SLICE_X141Y122_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X141Y122_AO6),
.Q(CLBLM_R_X89Y122_SLICE_X141Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X141Y122_BO6),
.Q(CLBLM_R_X89Y122_SLICE_X141Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y122_SLICE_X141Y122_DO6),
.Q(CLBLM_R_X89Y122_SLICE_X141Y122_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X89Y122_SLICE_X141Y122_BQ),
.I3(1'b1),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_DQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y122_SLICE_X141Y122_DO5),
.O6(CLBLM_R_X89Y122_SLICE_X141Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acc00cc00)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_CLUT (
.I0(CLBLM_R_X89Y122_SLICE_X141Y122_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X89Y122_SLICE_X141Y122_DQ),
.I3(CLBLM_R_X89Y121_SLICE_X141Y121_C5Q),
.I4(CLBLM_R_X89Y122_SLICE_X141Y122_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y122_SLICE_X141Y122_CO5),
.O6(CLBLM_R_X89Y122_SLICE_X141Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ee0000e4440000)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X92Y125_SLICE_X145Y125_DO6),
.I2(CLBLM_R_X89Y122_SLICE_X141Y122_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X89Y122_SLICE_X141Y122_CO6),
.O5(CLBLM_R_X89Y122_SLICE_X141Y122_BO5),
.O6(CLBLM_R_X89Y122_SLICE_X141Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X89Y122_SLICE_X141Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y124_SLICE_X141Y124_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y122_SLICE_X141Y122_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y122_SLICE_X141Y122_AO5),
.O6(CLBLM_R_X89Y122_SLICE_X141Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y123_SLICE_X140Y123_BO5),
.Q(CLBLM_R_X89Y123_SLICE_X140Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y123_SLICE_X140Y123_CO5),
.Q(CLBLM_R_X89Y123_SLICE_X140Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y123_SLICE_X140Y123_AO6),
.Q(CLBLM_R_X89Y123_SLICE_X140Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y123_SLICE_X140Y123_CO6),
.Q(CLBLM_R_X89Y123_SLICE_X140Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_DLUT (
.I0(CLBLM_R_X89Y123_SLICE_X140Y123_C5Q),
.I1(CLBLM_R_X89Y123_SLICE_X140Y123_AQ),
.I2(CLBLM_L_X92Y123_SLICE_X144Y123_D5Q),
.I3(CLBLM_R_X89Y123_SLICE_X140Y123_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y123_SLICE_X140Y123_CQ),
.O5(CLBLM_R_X89Y123_SLICE_X140Y123_DO5),
.O6(CLBLM_R_X89Y123_SLICE_X140Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y123_SLICE_X140Y123_CQ),
.I2(CLBLM_R_X89Y123_SLICE_X140Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y123_SLICE_X140Y123_CO5),
.O6(CLBLM_R_X89Y123_SLICE_X140Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_BLUT (
.I0(CLBLM_R_X89Y123_SLICE_X140Y123_AQ),
.I1(CLBLM_R_X89Y123_SLICE_X140Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y123_SLICE_X140Y123_CQ),
.I4(CLBLM_R_X89Y123_SLICE_X140Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y123_SLICE_X140Y123_BO5),
.O6(CLBLM_R_X89Y123_SLICE_X140Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaca00003a0a0000)
  ) CLBLM_R_X89Y123_SLICE_X140Y123_ALUT (
.I0(CLBLM_R_X89Y128_SLICE_X140Y128_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X89Y123_SLICE_X140Y123_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X89Y124_SLICE_X140Y124_A5Q),
.O5(CLBLM_R_X89Y123_SLICE_X140Y123_AO5),
.O6(CLBLM_R_X89Y123_SLICE_X140Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y123_SLICE_X141Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y123_SLICE_X141Y123_AO5),
.Q(CLBLM_R_X89Y123_SLICE_X141Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y123_SLICE_X141Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y123_SLICE_X141Y123_AO6),
.Q(CLBLM_R_X89Y123_SLICE_X141Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y123_SLICE_X141Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y123_SLICE_X141Y123_DO5),
.O6(CLBLM_R_X89Y123_SLICE_X141Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y123_SLICE_X141Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y123_SLICE_X141Y123_CO5),
.O6(CLBLM_R_X89Y123_SLICE_X141Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y123_SLICE_X141Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y123_SLICE_X141Y123_BO5),
.O6(CLBLM_R_X89Y123_SLICE_X141Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc030c030a0a05050)
  ) CLBLM_R_X89Y123_SLICE_X141Y123_ALUT (
.I0(CLBLM_R_X89Y123_SLICE_X141Y123_AQ),
.I1(CLBLM_L_X90Y121_SLICE_X143Y121_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y123_SLICE_X142Y123_BQ),
.I4(CLBLM_R_X89Y122_SLICE_X140Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y123_SLICE_X141Y123_AO5),
.O6(CLBLM_R_X89Y123_SLICE_X141Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X140Y124_AO5),
.Q(CLBLM_R_X89Y124_SLICE_X140Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X140Y124_AO6),
.Q(CLBLM_R_X89Y124_SLICE_X140Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X140Y124_BO5),
.Q(CLBLM_R_X89Y124_SLICE_X140Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X140Y124_CO6),
.Q(CLBLM_R_X89Y124_SLICE_X140Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5aa5cccca55a)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_DLUT (
.I0(CLBLM_R_X89Y122_SLICE_X141Y122_D5Q),
.I1(CLBLM_R_X89Y124_SLICE_X140Y124_CQ),
.I2(CLBLM_R_X89Y124_SLICE_X140Y124_BQ),
.I3(CLBLM_R_X89Y125_SLICE_X140Y125_DQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y124_SLICE_X141Y124_BQ),
.O5(CLBLM_R_X89Y124_SLICE_X140Y124_DO5),
.O6(CLBLM_R_X89Y124_SLICE_X140Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0000aaaa0000aa)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X89Y121_SLICE_X140Y121_A5Q),
.I4(CLBLM_R_X89Y126_SLICE_X140Y126_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y124_SLICE_X140Y124_CO5),
.O6(CLBLM_R_X89Y124_SLICE_X140Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_BLUT (
.I0(CLBLM_R_X89Y125_SLICE_X140Y125_DQ),
.I1(CLBLM_R_X89Y124_SLICE_X140Y124_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y124_SLICE_X141Y124_BQ),
.I4(CLBLM_R_X89Y122_SLICE_X141Y122_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y124_SLICE_X140Y124_BO5),
.O6(CLBLM_R_X89Y124_SLICE_X140Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0a0a0a0a0)
  ) CLBLM_R_X89Y124_SLICE_X140Y124_ALUT (
.I0(CLBLM_L_X90Y125_SLICE_X143Y125_AQ),
.I1(CLBLM_R_X89Y124_SLICE_X140Y124_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y124_SLICE_X140Y124_AO5),
.O6(CLBLM_R_X89Y124_SLICE_X140Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X141Y124_AO5),
.Q(CLBLM_R_X89Y124_SLICE_X141Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X141Y124_AO6),
.Q(CLBLM_R_X89Y124_SLICE_X141Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y124_SLICE_X141Y124_BO6),
.Q(CLBLM_R_X89Y124_SLICE_X141Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y124_SLICE_X141Y124_DO5),
.O6(CLBLM_R_X89Y124_SLICE_X141Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y124_SLICE_X141Y124_CO5),
.O6(CLBLM_R_X89Y124_SLICE_X141Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d050d0a0800080)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X89Y124_SLICE_X140Y124_BO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X89Y124_SLICE_X141Y124_A5Q),
.I5(CLBLM_L_X92Y127_SLICE_X145Y127_CO6),
.O5(CLBLM_R_X89Y124_SLICE_X141Y124_BO5),
.O6(CLBLM_R_X89Y124_SLICE_X141Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X89Y124_SLICE_X141Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y124_SLICE_X141Y124_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y130_SLICE_X141Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y124_SLICE_X141Y124_AO5),
.O6(CLBLM_R_X89Y124_SLICE_X141Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X140Y125_AO5),
.Q(CLBLM_R_X89Y125_SLICE_X140Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X140Y125_CO5),
.Q(CLBLM_R_X89Y125_SLICE_X140Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X140Y125_DO5),
.Q(CLBLM_R_X89Y125_SLICE_X140Y125_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X140Y125_AO6),
.Q(CLBLM_R_X89Y125_SLICE_X140Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X140Y125_BO6),
.Q(CLBLM_R_X89Y125_SLICE_X140Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X140Y125_DO6),
.Q(CLBLM_R_X89Y125_SLICE_X140Y125_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y128_SLICE_X140Y128_CQ),
.I2(CLBLM_R_X89Y124_SLICE_X141Y124_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y125_SLICE_X140Y125_DO5),
.O6(CLBLM_R_X89Y125_SLICE_X140Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caa00aa00)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X90Y125_SLICE_X142Y125_AQ),
.I2(CLBLM_R_X89Y125_SLICE_X140Y125_BQ),
.I3(CLBLM_R_X89Y125_SLICE_X141Y125_C5Q),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y125_SLICE_X140Y125_CO5),
.O6(CLBLM_R_X89Y125_SLICE_X140Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e020e0e0202020)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_BLUT (
.I0(CLBLM_R_X93Y126_SLICE_X147Y126_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_A5Q),
.I5(CLBLM_R_X89Y125_SLICE_X140Y125_CO6),
.O5(CLBLM_R_X89Y125_SLICE_X140Y125_BO5),
.O6(CLBLM_R_X89Y125_SLICE_X140Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c00000f0f0)
  ) CLBLM_R_X89Y125_SLICE_X140Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y125_SLICE_X140Y125_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_L_X90Y118_SLICE_X143Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y125_SLICE_X140Y125_AO5),
.O6(CLBLM_R_X89Y125_SLICE_X140Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X141Y125_BO5),
.Q(CLBLM_R_X89Y125_SLICE_X141Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X141Y125_CO5),
.Q(CLBLM_R_X89Y125_SLICE_X141Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X141Y125_AO6),
.Q(CLBLM_R_X89Y125_SLICE_X141Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y125_SLICE_X141Y125_CO6),
.Q(CLBLM_R_X89Y125_SLICE_X141Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_DLUT (
.I0(CLBLM_R_X89Y126_SLICE_X141Y126_C5Q),
.I1(CLBLM_R_X89Y125_SLICE_X141Y125_CQ),
.I2(CLBLM_R_X89Y125_SLICE_X141Y125_AQ),
.I3(CLBLM_R_X89Y125_SLICE_X141Y125_A5Q),
.I4(CLBLM_R_X89Y123_SLICE_X141Y123_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y125_SLICE_X141Y125_DO5),
.O6(CLBLM_R_X89Y125_SLICE_X141Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aa00aa00)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X90Y125_SLICE_X142Y125_AQ),
.I4(CLBLM_R_X89Y125_SLICE_X141Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y125_SLICE_X141Y125_CO5),
.O6(CLBLM_R_X89Y125_SLICE_X141Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_BLUT (
.I0(CLBLM_R_X89Y125_SLICE_X141Y125_AQ),
.I1(CLBLM_R_X89Y125_SLICE_X141Y125_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y125_SLICE_X141Y125_CQ),
.I4(CLBLM_R_X89Y126_SLICE_X141Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y125_SLICE_X141Y125_BO5),
.O6(CLBLM_R_X89Y125_SLICE_X141Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e04040e040e040)
  ) CLBLM_R_X89Y125_SLICE_X141Y125_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X92Y126_SLICE_X145Y126_DO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y125_SLICE_X141Y125_BO6),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X89Y125_SLICE_X141Y125_AO5),
.O6(CLBLM_R_X89Y125_SLICE_X141Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X140Y126_BO5),
.Q(CLBLM_R_X89Y126_SLICE_X140Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X140Y126_AO6),
.Q(CLBLM_R_X89Y126_SLICE_X140Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X140Y126_BO6),
.Q(CLBLM_R_X89Y126_SLICE_X140Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y126_SLICE_X140Y126_DO5),
.O6(CLBLM_R_X89Y126_SLICE_X140Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y126_SLICE_X140Y126_CO5),
.O6(CLBLM_R_X89Y126_SLICE_X140Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha050a050c0c03030)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_BLUT (
.I0(CLBLM_L_X90Y126_SLICE_X142Y126_AQ),
.I1(CLBLM_R_X89Y123_SLICE_X140Y123_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y126_SLICE_X142Y126_C5Q),
.I4(CLBLM_R_X89Y126_SLICE_X140Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y126_SLICE_X140Y126_BO5),
.O6(CLBLM_R_X89Y126_SLICE_X140Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0d050d0a0800080)
  ) CLBLM_R_X89Y126_SLICE_X140Y126_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_L_X90Y126_SLICE_X142Y126_AO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X90Y125_SLICE_X143Y125_AQ),
.I5(CLBLM_R_X89Y130_SLICE_X140Y130_BO6),
.O5(CLBLM_R_X89Y126_SLICE_X140Y126_AO5),
.O6(CLBLM_R_X89Y126_SLICE_X140Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X141Y126_BO5),
.Q(CLBLM_R_X89Y126_SLICE_X141Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X141Y126_CO5),
.Q(CLBLM_R_X89Y126_SLICE_X141Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X141Y126_AO6),
.Q(CLBLM_R_X89Y126_SLICE_X141Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y126_SLICE_X141Y126_CO6),
.Q(CLBLM_R_X89Y126_SLICE_X141Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_DLUT (
.I0(CLBLM_R_X89Y123_SLICE_X141Y123_A5Q),
.I1(CLBLM_R_X89Y128_SLICE_X141Y128_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X89Y126_SLICE_X141Y126_A5Q),
.I4(CLBLM_R_X89Y126_SLICE_X141Y126_AQ),
.I5(CLBLM_R_X89Y126_SLICE_X141Y126_CQ),
.O5(CLBLM_R_X89Y126_SLICE_X141Y126_DO5),
.O6(CLBLM_R_X89Y126_SLICE_X141Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X89Y125_SLICE_X141Y125_CQ),
.I3(1'b1),
.I4(CLBLM_R_X89Y126_SLICE_X141Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y126_SLICE_X141Y126_CO5),
.O6(CLBLM_R_X89Y126_SLICE_X141Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996aaaa0000)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_BLUT (
.I0(CLBLM_R_X89Y128_SLICE_X141Y128_A5Q),
.I1(CLBLM_R_X89Y126_SLICE_X141Y126_A5Q),
.I2(CLBLM_R_X89Y126_SLICE_X141Y126_AQ),
.I3(CLBLM_R_X89Y126_SLICE_X141Y126_CQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X89Y126_SLICE_X141Y126_BO5),
.O6(CLBLM_R_X89Y126_SLICE_X141Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b0c08070304000)
  ) CLBLM_R_X89Y126_SLICE_X141Y126_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y126_SLICE_X141Y126_BO6),
.I4(CLBLM_R_X93Y126_SLICE_X146Y126_DO6),
.I5(CLBLM_R_X89Y127_SLICE_X141Y127_A5Q),
.O5(CLBLM_R_X89Y126_SLICE_X141Y126_AO5),
.O6(CLBLM_R_X89Y126_SLICE_X141Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X140Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X140Y127_DO5),
.O6(CLBLM_R_X89Y127_SLICE_X140Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X140Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X140Y127_CO5),
.O6(CLBLM_R_X89Y127_SLICE_X140Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X140Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X140Y127_BO5),
.O6(CLBLM_R_X89Y127_SLICE_X140Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X140Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X140Y127_AO5),
.O6(CLBLM_R_X89Y127_SLICE_X140Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y127_SLICE_X141Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y127_SLICE_X141Y127_AO5),
.Q(CLBLM_R_X89Y127_SLICE_X141Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y127_SLICE_X141Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y127_SLICE_X141Y127_AO6),
.Q(CLBLM_R_X89Y127_SLICE_X141Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X141Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X141Y127_DO5),
.O6(CLBLM_R_X89Y127_SLICE_X141Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X141Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X141Y127_CO5),
.O6(CLBLM_R_X89Y127_SLICE_X141Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y127_SLICE_X141Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X141Y127_BO5),
.O6(CLBLM_R_X89Y127_SLICE_X141Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_R_X89Y127_SLICE_X141Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X89Y127_SLICE_X141Y127_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y127_SLICE_X141Y127_AO5),
.O6(CLBLM_R_X89Y127_SLICE_X141Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y128_SLICE_X140Y128_BO5),
.Q(CLBLM_R_X89Y128_SLICE_X140Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y128_SLICE_X140Y128_CO5),
.Q(CLBLM_R_X89Y128_SLICE_X140Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y128_SLICE_X140Y128_AO6),
.Q(CLBLM_R_X89Y128_SLICE_X140Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y128_SLICE_X140Y128_CO6),
.Q(CLBLM_R_X89Y128_SLICE_X140Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5aa5cccca55a)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_DLUT (
.I0(CLBLM_R_X89Y125_SLICE_X140Y125_D5Q),
.I1(CLBLM_R_X89Y126_SLICE_X140Y126_B5Q),
.I2(CLBLM_R_X89Y128_SLICE_X140Y128_AQ),
.I3(CLBLM_R_X89Y128_SLICE_X140Y128_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X89Y128_SLICE_X140Y128_CQ),
.O5(CLBLM_R_X89Y128_SLICE_X140Y128_DO5),
.O6(CLBLM_R_X89Y128_SLICE_X140Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y128_SLICE_X140Y128_AQ),
.I2(CLBLM_R_X89Y131_SLICE_X140Y131_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y128_SLICE_X140Y128_CO5),
.O6(CLBLM_R_X89Y128_SLICE_X140Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_BLUT (
.I0(CLBLM_R_X89Y128_SLICE_X140Y128_AQ),
.I1(CLBLM_R_X89Y128_SLICE_X140Y128_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y128_SLICE_X140Y128_CQ),
.I4(CLBLM_R_X89Y125_SLICE_X140Y125_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y128_SLICE_X140Y128_BO5),
.O6(CLBLM_R_X89Y128_SLICE_X140Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c03000a0a0a0a0)
  ) CLBLM_R_X89Y128_SLICE_X140Y128_ALUT (
.I0(CLBLM_R_X93Y130_SLICE_X147Y130_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y128_SLICE_X140Y128_BO6),
.I4(CLBLM_R_X89Y130_SLICE_X141Y130_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X89Y128_SLICE_X140Y128_AO5),
.O6(CLBLM_R_X89Y128_SLICE_X140Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y128_SLICE_X141Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y128_SLICE_X141Y128_AO5),
.Q(CLBLM_R_X89Y128_SLICE_X141Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y128_SLICE_X141Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y128_SLICE_X141Y128_AO6),
.Q(CLBLM_R_X89Y128_SLICE_X141Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y128_SLICE_X141Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y128_SLICE_X141Y128_DO5),
.O6(CLBLM_R_X89Y128_SLICE_X141Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y128_SLICE_X141Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y128_SLICE_X141Y128_CO5),
.O6(CLBLM_R_X89Y128_SLICE_X141Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y128_SLICE_X141Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y128_SLICE_X141Y128_BO5),
.O6(CLBLM_R_X89Y128_SLICE_X141Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f000f000)
  ) CLBLM_R_X89Y128_SLICE_X141Y128_ALUT (
.I0(CLBLM_L_X90Y128_SLICE_X143Y128_CQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X89Y126_SLICE_X141Y126_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y128_SLICE_X141Y128_AO5),
.O6(CLBLM_R_X89Y128_SLICE_X141Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y130_SLICE_X140Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y130_SLICE_X140Y130_AO5),
.Q(CLBLM_R_X89Y130_SLICE_X140Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y130_SLICE_X140Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y130_SLICE_X140Y130_DO5),
.O6(CLBLM_R_X89Y130_SLICE_X140Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y130_SLICE_X140Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y130_SLICE_X140Y130_CO5),
.O6(CLBLM_R_X89Y130_SLICE_X140Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X89Y130_SLICE_X140Y130_BLUT (
.I0(CLBLM_R_X89Y131_SLICE_X140Y131_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X89Y130_SLICE_X140Y130_AQ),
.I3(CLBLM_R_X89Y130_SLICE_X141Y130_BQ),
.I4(CLBLM_R_X89Y128_SLICE_X140Y128_C5Q),
.I5(CLBLM_R_X89Y126_SLICE_X140Y126_BQ),
.O5(CLBLM_R_X89Y130_SLICE_X140Y130_BO5),
.O6(CLBLM_R_X89Y130_SLICE_X140Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_R_X89Y130_SLICE_X140Y130_ALUT (
.I0(CLBLM_R_X89Y130_SLICE_X141Y130_BQ),
.I1(CLBLM_R_X89Y131_SLICE_X140Y131_AQ),
.I2(CLBLM_R_X89Y130_SLICE_X140Y130_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X89Y128_SLICE_X140Y128_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X89Y130_SLICE_X140Y130_AO5),
.O6(CLBLM_R_X89Y130_SLICE_X140Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y130_SLICE_X141Y130_AO5),
.Q(CLBLM_R_X89Y130_SLICE_X141Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y130_SLICE_X141Y130_AO6),
.Q(CLBLM_R_X89Y130_SLICE_X141Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y130_SLICE_X141Y130_BO6),
.Q(CLBLM_R_X89Y130_SLICE_X141Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y130_SLICE_X141Y130_DO5),
.O6(CLBLM_R_X89Y130_SLICE_X141Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y130_SLICE_X141Y130_CO5),
.O6(CLBLM_R_X89Y130_SLICE_X141Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaf0aa00000000)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_BLUT (
.I0(CLBLM_L_X92Y132_SLICE_X145Y132_DO6),
.I1(CLBLM_R_X89Y130_SLICE_X141Y130_A5Q),
.I2(CLBLM_R_X89Y130_SLICE_X140Y130_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X89Y130_SLICE_X141Y130_BO5),
.O6(CLBLM_R_X89Y130_SLICE_X141Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X89Y130_SLICE_X141Y130_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X89Y130_SLICE_X141Y130_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X90Y130_SLICE_X142Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y130_SLICE_X141Y130_AO5),
.O6(CLBLM_R_X89Y130_SLICE_X141Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y131_SLICE_X140Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y131_SLICE_X140Y131_AO5),
.Q(CLBLM_R_X89Y131_SLICE_X140Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X89Y131_SLICE_X140Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X89Y131_SLICE_X140Y131_AO6),
.Q(CLBLM_R_X89Y131_SLICE_X140Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X140Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X140Y131_DO5),
.O6(CLBLM_R_X89Y131_SLICE_X140Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X140Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X140Y131_CO5),
.O6(CLBLM_R_X89Y131_SLICE_X140Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X140Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X140Y131_BO5),
.O6(CLBLM_R_X89Y131_SLICE_X140Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000aa00aa00)
  ) CLBLM_R_X89Y131_SLICE_X140Y131_ALUT (
.I0(CLBLM_L_X90Y131_SLICE_X142Y131_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X89Y130_SLICE_X141Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X140Y131_AO5),
.O6(CLBLM_R_X89Y131_SLICE_X140Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X141Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X141Y131_DO5),
.O6(CLBLM_R_X89Y131_SLICE_X141Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X141Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X141Y131_CO5),
.O6(CLBLM_R_X89Y131_SLICE_X141Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X141Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X141Y131_BO5),
.O6(CLBLM_R_X89Y131_SLICE_X141Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X89Y131_SLICE_X141Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X89Y131_SLICE_X141Y131_AO5),
.O6(CLBLM_R_X89Y131_SLICE_X141Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y111_SLICE_X146Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X146Y111_DO5),
.O6(CLBLM_R_X93Y111_SLICE_X146Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y111_SLICE_X146Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X146Y111_CO5),
.O6(CLBLM_R_X93Y111_SLICE_X146Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y111_SLICE_X146Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X146Y111_BO5),
.O6(CLBLM_R_X93Y111_SLICE_X146Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y111_SLICE_X146Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X146Y111_AO5),
.O6(CLBLM_R_X93Y111_SLICE_X146Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y111_SLICE_X147Y111_AO5),
.Q(CLBLM_R_X93Y111_SLICE_X147Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y111_SLICE_X147Y111_BO5),
.Q(CLBLM_R_X93Y111_SLICE_X147Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y111_SLICE_X147Y111_AO6),
.Q(CLBLM_R_X93Y111_SLICE_X147Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y111_SLICE_X147Y111_BO6),
.Q(CLBLM_R_X93Y111_SLICE_X147Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X147Y111_DO5),
.O6(CLBLM_R_X93Y111_SLICE_X147Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y111_SLICE_X147Y111_AQ),
.I2(CLBLM_R_X93Y111_SLICE_X147Y111_BQ),
.I3(CLBLM_R_X93Y112_SLICE_X147Y112_BQ),
.I4(CLBLM_R_X93Y111_SLICE_X147Y111_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X147Y111_CO5),
.O6(CLBLM_R_X93Y111_SLICE_X147Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y111_SLICE_X147Y111_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y111_SLICE_X147Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X147Y111_BO5),
.O6(CLBLM_R_X93Y111_SLICE_X147Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_R_X93Y111_SLICE_X147Y111_ALUT (
.I0(CLBLM_R_X93Y112_SLICE_X147Y112_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y112_SLICE_X146Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y111_SLICE_X147Y111_AO5),
.O6(CLBLM_R_X93Y111_SLICE_X147Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X146Y112_AO5),
.Q(CLBLM_R_X93Y112_SLICE_X146Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X146Y112_BO5),
.Q(CLBLM_R_X93Y112_SLICE_X146Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X146Y112_AO6),
.Q(CLBLM_R_X93Y112_SLICE_X146Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X146Y112_BO6),
.Q(CLBLM_R_X93Y112_SLICE_X146Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_L_X92Y112_SLICE_X145Y112_A5Q),
.I3(CLBLM_R_X93Y112_SLICE_X146Y112_BQ),
.I4(CLBLM_R_X93Y112_SLICE_X146Y112_B5Q),
.I5(CLBLM_R_X93Y115_SLICE_X146Y115_BQ),
.O5(CLBLM_R_X93Y112_SLICE_X146Y112_DO5),
.O6(CLBLM_R_X93Y112_SLICE_X146Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y111_SLICE_X147Y111_A5Q),
.I2(CLBLM_R_X93Y112_SLICE_X146Y112_AQ),
.I3(CLBLM_R_X93Y112_SLICE_X146Y112_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X94Y112_SLICE_X148Y112_BQ),
.O5(CLBLM_R_X93Y112_SLICE_X146Y112_CO5),
.O6(CLBLM_R_X93Y112_SLICE_X146Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_BLUT (
.I0(CLBLM_R_X93Y112_SLICE_X146Y112_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y115_SLICE_X146Y115_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y112_SLICE_X146Y112_BO5),
.O6(CLBLM_R_X93Y112_SLICE_X146Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X93Y112_SLICE_X146Y112_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y112_SLICE_X146Y112_AQ),
.I3(1'b1),
.I4(CLBLM_L_X94Y112_SLICE_X148Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y112_SLICE_X146Y112_AO5),
.O6(CLBLM_R_X93Y112_SLICE_X146Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X147Y112_AO5),
.Q(CLBLM_R_X93Y112_SLICE_X147Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X147Y112_BO5),
.Q(CLBLM_R_X93Y112_SLICE_X147Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X147Y112_CO5),
.Q(CLBLM_R_X93Y112_SLICE_X147Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X147Y112_AO6),
.Q(CLBLM_R_X93Y112_SLICE_X147Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X147Y112_BO6),
.Q(CLBLM_R_X93Y112_SLICE_X147Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y112_SLICE_X147Y112_CO6),
.Q(CLBLM_R_X93Y112_SLICE_X147Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_DLUT (
.I0(CLBLM_R_X93Y112_SLICE_X147Y112_C5Q),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_CQ),
.I2(1'b1),
.I3(CLBLM_R_X93Y114_SLICE_X147Y114_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X94Y115_SLICE_X148Y115_CQ),
.O5(CLBLM_R_X93Y112_SLICE_X147Y112_DO5),
.O6(CLBLM_R_X93Y112_SLICE_X147Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_CQ),
.I2(1'b1),
.I3(CLBLM_R_X93Y114_SLICE_X147Y114_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y112_SLICE_X147Y112_CO5),
.O6(CLBLM_R_X93Y112_SLICE_X147Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0000a5a50000)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_BLUT (
.I0(CLBLM_L_X94Y112_SLICE_X148Y112_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X93Y113_SLICE_X147Y113_B5Q),
.I3(CLBLM_L_X94Y112_SLICE_X148Y112_CO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X93Y112_SLICE_X147Y112_BO5),
.O6(CLBLM_R_X93Y112_SLICE_X147Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X93Y112_SLICE_X147Y112_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y112_SLICE_X148Y112_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y112_SLICE_X147Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y112_SLICE_X147Y112_AO5),
.O6(CLBLM_R_X93Y112_SLICE_X147Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X146Y113_AO5),
.Q(CLBLM_R_X93Y113_SLICE_X146Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X146Y113_BO5),
.Q(CLBLM_R_X93Y113_SLICE_X146Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X146Y113_AO6),
.Q(CLBLM_R_X93Y113_SLICE_X146Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X146Y113_BO6),
.Q(CLBLM_R_X93Y113_SLICE_X146Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y113_SLICE_X146Y113_AQ),
.I2(CLBLM_L_X92Y113_SLICE_X144Y113_A5Q),
.I3(CLBLM_R_X93Y113_SLICE_X146Y113_BQ),
.I4(CLBLM_R_X93Y113_SLICE_X146Y113_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y113_SLICE_X146Y113_DO5),
.O6(CLBLM_R_X93Y113_SLICE_X146Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03cf03cfeeee2222)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_CLUT (
.I0(CLBLM_L_X92Y112_SLICE_X145Y112_CO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X94Y113_SLICE_X148Y113_A5Q),
.I3(CLBLM_R_X93Y112_SLICE_X147Y112_A5Q),
.I4(CLBLM_R_X93Y113_SLICE_X146Y113_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X93Y113_SLICE_X146Y113_CO5),
.O6(CLBLM_R_X93Y113_SLICE_X146Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y113_SLICE_X146Y113_BQ),
.I2(CLBLM_R_X93Y113_SLICE_X146Y113_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y113_SLICE_X146Y113_BO5),
.O6(CLBLM_R_X93Y113_SLICE_X146Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330000aa550000)
  ) CLBLM_R_X93Y113_SLICE_X146Y113_ALUT (
.I0(CLBLM_L_X92Y112_SLICE_X145Y112_A5Q),
.I1(CLBLM_R_X93Y113_SLICE_X146Y113_CO6),
.I2(1'b1),
.I3(CLBLM_R_X93Y112_SLICE_X147Y112_B5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X93Y113_SLICE_X146Y113_AO5),
.O6(CLBLM_R_X93Y113_SLICE_X146Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X147Y113_AO5),
.Q(CLBLM_R_X93Y113_SLICE_X147Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X147Y113_BO5),
.Q(CLBLM_R_X93Y113_SLICE_X147Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X147Y113_AO6),
.Q(CLBLM_R_X93Y113_SLICE_X147Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y113_SLICE_X147Y113_BO6),
.Q(CLBLM_R_X93Y113_SLICE_X147Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y113_SLICE_X147Y113_AQ),
.I2(CLBLM_R_X93Y113_SLICE_X147Y113_BQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y113_SLICE_X147Y113_B5Q),
.I5(CLBLM_R_X93Y115_SLICE_X147Y115_BQ),
.O5(CLBLM_R_X93Y113_SLICE_X147Y113_DO5),
.O6(CLBLM_R_X93Y113_SLICE_X147Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h53535353fff00f00)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_CLUT (
.I0(CLBLM_L_X94Y113_SLICE_X148Y113_BQ),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_B5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y119_SLICE_X149Y119_DO6),
.I4(CLBLM_R_X93Y113_SLICE_X147Y113_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X93Y113_SLICE_X147Y113_CO5),
.O6(CLBLM_R_X93Y113_SLICE_X147Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y113_SLICE_X147Y113_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y113_SLICE_X147Y113_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y113_SLICE_X147Y113_BO5),
.O6(CLBLM_R_X93Y113_SLICE_X147Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X93Y113_SLICE_X147Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y115_SLICE_X147Y115_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X94Y114_SLICE_X148Y114_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y113_SLICE_X147Y113_AO5),
.O6(CLBLM_R_X93Y113_SLICE_X147Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X146Y114_AO5),
.Q(CLBLM_R_X93Y114_SLICE_X146Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X146Y114_BO5),
.Q(CLBLM_R_X93Y114_SLICE_X146Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X146Y114_AO6),
.Q(CLBLM_R_X93Y114_SLICE_X146Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X146Y114_BO6),
.Q(CLBLM_R_X93Y114_SLICE_X146Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0cfa0c0afcfafc)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_DLUT (
.I0(CLBLM_L_X90Y113_SLICE_X143Y113_DO6),
.I1(CLBLM_R_X93Y116_SLICE_X147Y116_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X92Y114_SLICE_X145Y114_A5Q),
.I5(CLBLM_L_X90Y113_SLICE_X143Y113_A5Q),
.O5(CLBLM_R_X93Y114_SLICE_X146Y114_DO5),
.O6(CLBLM_R_X93Y114_SLICE_X146Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f303f300a0afafa)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_CLUT (
.I0(CLBLM_L_X90Y113_SLICE_X143Y113_DO6),
.I1(CLBLM_R_X93Y112_SLICE_X147Y112_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X92Y113_SLICE_X144Y113_CO6),
.I4(CLBLM_R_X93Y115_SLICE_X147Y115_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X93Y114_SLICE_X146Y114_CO5),
.O6(CLBLM_R_X93Y114_SLICE_X146Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f090909090)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_BLUT (
.I0(CLBLM_R_X93Y115_SLICE_X146Y115_A5Q),
.I1(CLBLM_R_X93Y116_SLICE_X147Y116_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y114_SLICE_X146Y114_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y114_SLICE_X146Y114_BO5),
.O6(CLBLM_R_X93Y114_SLICE_X146Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030a050a050)
  ) CLBLM_R_X93Y114_SLICE_X146Y114_ALUT (
.I0(CLBLM_R_X93Y116_SLICE_X147Y116_B5Q),
.I1(CLBLM_L_X92Y114_SLICE_X144Y114_CO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y114_SLICE_X146Y114_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y114_SLICE_X146Y114_AO5),
.O6(CLBLM_R_X93Y114_SLICE_X146Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X147Y114_AO5),
.Q(CLBLM_R_X93Y114_SLICE_X147Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X147Y114_BO5),
.Q(CLBLM_R_X93Y114_SLICE_X147Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X147Y114_AO6),
.Q(CLBLM_R_X93Y114_SLICE_X147Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y114_SLICE_X147Y114_BO6),
.Q(CLBLM_R_X93Y114_SLICE_X147Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y114_SLICE_X147Y114_DO5),
.O6(CLBLM_R_X93Y114_SLICE_X147Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_R_X93Y114_SLICE_X147Y114_BQ),
.I3(CLBLM_R_X93Y114_SLICE_X147Y114_A5Q),
.I4(CLBLM_R_X93Y114_SLICE_X147Y114_B5Q),
.I5(CLBLM_L_X94Y115_SLICE_X149Y115_AQ),
.O5(CLBLM_R_X93Y114_SLICE_X147Y114_CO5),
.O6(CLBLM_R_X93Y114_SLICE_X147Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y114_SLICE_X147Y114_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X94Y115_SLICE_X149Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y114_SLICE_X147Y114_BO5),
.O6(CLBLM_R_X93Y114_SLICE_X147Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X93Y114_SLICE_X147Y114_ALUT (
.I0(CLBLM_R_X93Y114_SLICE_X147Y114_B5Q),
.I1(CLBLM_L_X94Y115_SLICE_X148Y115_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y114_SLICE_X147Y114_AO5),
.O6(CLBLM_R_X93Y114_SLICE_X147Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X146Y115_AO5),
.Q(CLBLM_R_X93Y115_SLICE_X146Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X146Y115_BO5),
.Q(CLBLM_R_X93Y115_SLICE_X146Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X146Y115_AO6),
.Q(CLBLM_R_X93Y115_SLICE_X146Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X146Y115_BO6),
.Q(CLBLM_R_X93Y115_SLICE_X146Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X146Y115_DO5),
.O6(CLBLM_R_X93Y115_SLICE_X146Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X146Y115_CO5),
.O6(CLBLM_R_X93Y115_SLICE_X146Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc84848484)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_BLUT (
.I0(CLBLM_R_X93Y118_SLICE_X147Y118_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y115_SLICE_X147Y115_B5Q),
.I3(CLBLM_L_X92Y113_SLICE_X145Y113_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X146Y115_BO5),
.O6(CLBLM_R_X93Y115_SLICE_X146Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300a500a500)
  ) CLBLM_R_X93Y115_SLICE_X146Y115_ALUT (
.I0(CLBLM_R_X93Y115_SLICE_X146Y115_B5Q),
.I1(CLBLM_L_X92Y113_SLICE_X145Y113_CO6),
.I2(CLBLM_R_X93Y118_SLICE_X147Y118_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X146Y115_AO5),
.O6(CLBLM_R_X93Y115_SLICE_X146Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X147Y115_AO5),
.Q(CLBLM_R_X93Y115_SLICE_X147Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X147Y115_BO5),
.Q(CLBLM_R_X93Y115_SLICE_X147Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X147Y115_AO6),
.Q(CLBLM_R_X93Y115_SLICE_X147Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y115_SLICE_X147Y115_BO6),
.Q(CLBLM_R_X93Y115_SLICE_X147Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X147Y115_DO5),
.O6(CLBLM_R_X93Y115_SLICE_X147Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5404f4a45e0efeae)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X90Y113_SLICE_X142Y113_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X94Y115_SLICE_X148Y115_DO6),
.I4(CLBLM_L_X94Y114_SLICE_X149Y114_AQ),
.I5(CLBLM_R_X97Y115_SLICE_X152Y115_A5Q),
.O5(CLBLM_R_X93Y115_SLICE_X147Y115_CO5),
.O6(CLBLM_R_X93Y115_SLICE_X147Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00c300c300)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y116_SLICE_X148Y116_B5Q),
.I2(CLBLM_L_X94Y115_SLICE_X148Y115_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y113_SLICE_X147Y113_CO6),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X147Y115_BO5),
.O6(CLBLM_R_X93Y115_SLICE_X147Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00a500a500)
  ) CLBLM_R_X93Y115_SLICE_X147Y115_ALUT (
.I0(CLBLM_L_X94Y113_SLICE_X148Y113_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X92Y113_SLICE_X144Y113_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y115_SLICE_X147Y115_CO6),
.I5(1'b1),
.O5(CLBLM_R_X93Y115_SLICE_X147Y115_AO5),
.O6(CLBLM_R_X93Y115_SLICE_X147Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X146Y116_AO5),
.Q(CLBLM_R_X93Y116_SLICE_X146Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X146Y116_BO5),
.Q(CLBLM_R_X93Y116_SLICE_X146Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X146Y116_AO6),
.Q(CLBLM_R_X93Y116_SLICE_X146Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X146Y116_BO6),
.Q(CLBLM_R_X93Y116_SLICE_X146Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_DO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_CLUT (
.I0(CLBLM_L_X92Y115_SLICE_X145Y115_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X93Y116_SLICE_X146Y116_BQ),
.I3(CLBLM_R_X93Y116_SLICE_X146Y116_A5Q),
.I4(CLBLM_R_X93Y116_SLICE_X146Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_CO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_BLUT (
.I0(CLBLM_R_X93Y116_SLICE_X146Y116_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X92Y115_SLICE_X145Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_BO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X93Y116_SLICE_X146Y116_ALUT (
.I0(CLBLM_R_X93Y116_SLICE_X146Y116_B5Q),
.I1(CLBLM_L_X90Y115_SLICE_X143Y115_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X146Y116_AO5),
.O6(CLBLM_R_X93Y116_SLICE_X146Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X147Y116_AO5),
.Q(CLBLM_R_X93Y116_SLICE_X147Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X147Y116_BO5),
.Q(CLBLM_R_X93Y116_SLICE_X147Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X147Y116_AO6),
.Q(CLBLM_R_X93Y116_SLICE_X147Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y116_SLICE_X147Y116_BO6),
.Q(CLBLM_R_X93Y116_SLICE_X147Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_DO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_CLUT (
.I0(CLBLM_R_X93Y116_SLICE_X147Y116_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y116_SLICE_X147Y116_AQ),
.I4(CLBLM_R_X93Y116_SLICE_X147Y116_B5Q),
.I5(CLBLM_L_X94Y120_SLICE_X149Y120_AQ),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_CO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y116_SLICE_X147Y116_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y116_SLICE_X147Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_BO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X93Y116_SLICE_X147Y116_ALUT (
.I0(CLBLM_L_X94Y116_SLICE_X148Y116_A5Q),
.I1(CLBLM_L_X94Y120_SLICE_X149Y120_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y116_SLICE_X147Y116_AO5),
.O6(CLBLM_R_X93Y116_SLICE_X147Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y117_SLICE_X146Y117_AO5),
.Q(CLBLM_R_X93Y117_SLICE_X146Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y117_SLICE_X146Y117_BO5),
.Q(CLBLM_R_X93Y117_SLICE_X146Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y117_SLICE_X146Y117_AO6),
.Q(CLBLM_R_X93Y117_SLICE_X146Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y117_SLICE_X146Y117_BO6),
.Q(CLBLM_R_X93Y117_SLICE_X146Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X146Y117_DO5),
.O6(CLBLM_R_X93Y117_SLICE_X146Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_CLUT (
.I0(CLBLM_R_X93Y116_SLICE_X146Y116_AQ),
.I1(1'b1),
.I2(CLBLM_R_X93Y117_SLICE_X146Y117_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X93Y117_SLICE_X146Y117_B5Q),
.I5(CLBLM_L_X90Y115_SLICE_X143Y115_BQ),
.O5(CLBLM_R_X93Y117_SLICE_X146Y117_CO5),
.O6(CLBLM_R_X93Y117_SLICE_X146Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y117_SLICE_X146Y117_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y116_SLICE_X146Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X146Y117_BO5),
.O6(CLBLM_R_X93Y117_SLICE_X146Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88228822)
  ) CLBLM_R_X93Y117_SLICE_X146Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y117_SLICE_X146Y117_B5Q),
.I2(CLBLM_R_X97Y117_SLICE_X152Y117_CO6),
.I3(CLBLM_L_X94Y116_SLICE_X149Y116_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X146Y117_AO5),
.O6(CLBLM_R_X93Y117_SLICE_X146Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y117_SLICE_X147Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X147Y117_DO5),
.O6(CLBLM_R_X93Y117_SLICE_X147Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y117_SLICE_X147Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X147Y117_CO5),
.O6(CLBLM_R_X93Y117_SLICE_X147Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y117_SLICE_X147Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X147Y117_BO5),
.O6(CLBLM_R_X93Y117_SLICE_X147Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y117_SLICE_X147Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y117_SLICE_X147Y117_AO5),
.O6(CLBLM_R_X93Y117_SLICE_X147Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y118_SLICE_X146Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X146Y118_DO5),
.O6(CLBLM_R_X93Y118_SLICE_X146Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y118_SLICE_X146Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X146Y118_CO5),
.O6(CLBLM_R_X93Y118_SLICE_X146Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y118_SLICE_X146Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X146Y118_BO5),
.O6(CLBLM_R_X93Y118_SLICE_X146Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y118_SLICE_X146Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X146Y118_AO5),
.O6(CLBLM_R_X93Y118_SLICE_X146Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y118_SLICE_X147Y118_AO5),
.Q(CLBLM_R_X93Y118_SLICE_X147Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y118_SLICE_X147Y118_BO5),
.Q(CLBLM_R_X93Y118_SLICE_X147Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y118_SLICE_X147Y118_AO6),
.Q(CLBLM_R_X93Y118_SLICE_X147Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y118_SLICE_X147Y118_BO6),
.Q(CLBLM_R_X93Y118_SLICE_X147Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X147Y118_DO5),
.O6(CLBLM_R_X93Y118_SLICE_X147Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_CLUT (
.I0(CLBLM_L_X94Y119_SLICE_X149Y119_AQ),
.I1(CLBLM_R_X93Y118_SLICE_X147Y118_AQ),
.I2(CLBLM_R_X93Y118_SLICE_X147Y118_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X93Y118_SLICE_X147Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X147Y118_CO5),
.O6(CLBLM_R_X93Y118_SLICE_X147Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y118_SLICE_X147Y118_BQ),
.I2(CLBLM_R_X93Y118_SLICE_X147Y118_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X147Y118_BO5),
.O6(CLBLM_R_X93Y118_SLICE_X147Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X93Y118_SLICE_X147Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y119_SLICE_X149Y119_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X94Y119_SLICE_X149Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y118_SLICE_X147Y118_AO5),
.O6(CLBLM_R_X93Y118_SLICE_X147Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X146Y119_AO5),
.Q(CLBLM_R_X93Y119_SLICE_X146Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X146Y119_BO5),
.Q(CLBLM_R_X93Y119_SLICE_X146Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X146Y119_CO5),
.Q(CLBLM_R_X93Y119_SLICE_X146Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X146Y119_AO6),
.Q(CLBLM_R_X93Y119_SLICE_X146Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X146Y119_BO6),
.Q(CLBLM_R_X93Y119_SLICE_X146Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X146Y119_CO6),
.Q(CLBLM_R_X93Y119_SLICE_X146Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_DLUT (
.I0(CLBLM_R_X93Y119_SLICE_X146Y119_C5Q),
.I1(CLBLM_R_X93Y119_SLICE_X146Y119_CQ),
.I2(CLBLM_R_X93Y119_SLICE_X147Y119_AQ),
.I3(1'b1),
.I4(CLBLM_L_X94Y122_SLICE_X149Y122_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X93Y119_SLICE_X146Y119_DO5),
.O6(CLBLM_R_X93Y119_SLICE_X146Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_CLUT (
.I0(CLBLM_R_X93Y119_SLICE_X147Y119_AQ),
.I1(CLBLM_R_X93Y119_SLICE_X146Y119_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y119_SLICE_X146Y119_CO5),
.O6(CLBLM_R_X93Y119_SLICE_X146Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y114_SLICE_X146Y114_A5Q),
.I2(CLBLM_R_X93Y119_SLICE_X147Y119_A5Q),
.I3(CLBLM_L_X90Y118_SLICE_X143Y118_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y119_SLICE_X146Y119_BO5),
.O6(CLBLM_R_X93Y119_SLICE_X146Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0aaa0000aa)
  ) CLBLM_R_X93Y119_SLICE_X146Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X90Y119_SLICE_X143Y119_DO6),
.I3(CLBLM_R_X93Y119_SLICE_X146Y119_B5Q),
.I4(CLBLM_R_X93Y119_SLICE_X146Y119_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y119_SLICE_X146Y119_AO5),
.O6(CLBLM_R_X93Y119_SLICE_X146Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X147Y119_AO5),
.Q(CLBLM_R_X93Y119_SLICE_X147Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X147Y119_BO5),
.Q(CLBLM_R_X93Y119_SLICE_X147Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X147Y119_AO6),
.Q(CLBLM_R_X93Y119_SLICE_X147Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y119_SLICE_X147Y119_BO6),
.Q(CLBLM_R_X93Y119_SLICE_X147Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y119_SLICE_X147Y119_DO5),
.O6(CLBLM_R_X93Y119_SLICE_X147Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_CLUT (
.I0(CLBLM_R_X93Y119_SLICE_X147Y119_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y119_SLICE_X147Y119_A5Q),
.I4(CLBLM_R_X93Y119_SLICE_X147Y119_B5Q),
.I5(CLBLM_L_X94Y122_SLICE_X149Y122_BQ),
.O5(CLBLM_R_X93Y119_SLICE_X147Y119_CO5),
.O6(CLBLM_R_X93Y119_SLICE_X147Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaaa0000)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X94Y122_SLICE_X149Y122_BQ),
.I4(CLBLM_R_X93Y119_SLICE_X147Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y119_SLICE_X147Y119_BO5),
.O6(CLBLM_R_X93Y119_SLICE_X147Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aa00aa00)
  ) CLBLM_R_X93Y119_SLICE_X147Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X93Y119_SLICE_X147Y119_B5Q),
.I4(CLBLM_L_X94Y122_SLICE_X149Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y119_SLICE_X147Y119_AO5),
.O6(CLBLM_R_X93Y119_SLICE_X147Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X146Y120_AO5),
.Q(CLBLM_R_X93Y120_SLICE_X146Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X146Y120_BO5),
.Q(CLBLM_R_X93Y120_SLICE_X146Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X146Y120_AO6),
.Q(CLBLM_R_X93Y120_SLICE_X146Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X146Y120_BO6),
.Q(CLBLM_R_X93Y120_SLICE_X146Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X93Y120_SLICE_X147Y120_A5Q),
.I2(CLBLM_R_X93Y120_SLICE_X146Y120_BQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y120_SLICE_X146Y120_B5Q),
.I5(CLBLM_L_X94Y120_SLICE_X148Y120_CQ),
.O5(CLBLM_R_X93Y120_SLICE_X146Y120_DO5),
.O6(CLBLM_R_X93Y120_SLICE_X146Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05cf05c0f5cff5c0)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_CLUT (
.I0(CLBLM_L_X92Y119_SLICE_X144Y119_C5Q),
.I1(CLBLM_L_X92Y119_SLICE_X145Y119_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X95Y122_SLICE_X150Y122_DO6),
.I5(CLBLM_L_X92Y120_SLICE_X144Y120_AQ),
.O5(CLBLM_R_X93Y120_SLICE_X146Y120_CO5),
.O6(CLBLM_R_X93Y120_SLICE_X146Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y120_SLICE_X146Y120_BQ),
.I2(1'b1),
.I3(CLBLM_L_X94Y120_SLICE_X148Y120_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y120_SLICE_X146Y120_BO5),
.O6(CLBLM_R_X93Y120_SLICE_X146Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaa0a00a0a)
  ) CLBLM_R_X93Y120_SLICE_X146Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X93Y119_SLICE_X146Y119_A5Q),
.I3(CLBLM_L_X92Y120_SLICE_X144Y120_CO6),
.I4(CLBLM_R_X93Y124_SLICE_X147Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y120_SLICE_X146Y120_AO5),
.O6(CLBLM_R_X93Y120_SLICE_X146Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X147Y120_AO5),
.Q(CLBLM_R_X93Y120_SLICE_X147Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X147Y120_BO5),
.Q(CLBLM_R_X93Y120_SLICE_X147Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X147Y120_CO5),
.Q(CLBLM_R_X93Y120_SLICE_X147Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X147Y120_AO6),
.Q(CLBLM_R_X93Y120_SLICE_X147Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X147Y120_BO6),
.Q(CLBLM_R_X93Y120_SLICE_X147Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y120_SLICE_X147Y120_CO6),
.Q(CLBLM_R_X93Y120_SLICE_X147Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_DLUT (
.I0(CLBLM_L_X94Y120_SLICE_X148Y120_BQ),
.I1(1'b1),
.I2(CLBLM_R_X93Y120_SLICE_X147Y120_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X93Y120_SLICE_X147Y120_B5Q),
.I5(CLBLM_R_X93Y120_SLICE_X147Y120_AQ),
.O5(CLBLM_R_X93Y120_SLICE_X147Y120_DO5),
.O6(CLBLM_R_X93Y120_SLICE_X147Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha500a500cc003300)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_CLUT (
.I0(CLBLM_R_X93Y120_SLICE_X147Y120_A5Q),
.I1(CLBLM_R_X93Y120_SLICE_X147Y120_CQ),
.I2(CLBLM_L_X92Y119_SLICE_X144Y119_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y120_SLICE_X147Y120_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y120_SLICE_X147Y120_CO5),
.O6(CLBLM_R_X93Y120_SLICE_X147Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y120_SLICE_X147Y120_BQ),
.I2(CLBLM_R_X93Y120_SLICE_X147Y120_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y120_SLICE_X147Y120_BO5),
.O6(CLBLM_R_X93Y120_SLICE_X147Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaaa0000)
  ) CLBLM_R_X93Y120_SLICE_X147Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X94Y120_SLICE_X148Y120_BQ),
.I4(CLBLM_R_X93Y120_SLICE_X146Y120_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y120_SLICE_X147Y120_AO5),
.O6(CLBLM_R_X93Y120_SLICE_X147Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X146Y121_AO5),
.Q(CLBLM_R_X93Y121_SLICE_X146Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X146Y121_AO6),
.Q(CLBLM_R_X93Y121_SLICE_X146Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X146Y121_BO5),
.Q(CLBLM_R_X93Y121_SLICE_X146Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X146Y121_CO6),
.Q(CLBLM_R_X93Y121_SLICE_X146Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff690069ff960096)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_DLUT (
.I0(CLBLM_L_X92Y121_SLICE_X144Y121_BQ),
.I1(CLBLM_R_X93Y122_SLICE_X147Y122_C5Q),
.I2(CLBLM_R_X93Y121_SLICE_X146Y121_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y121_SLICE_X153Y121_CQ),
.I5(CLBLM_R_X93Y121_SLICE_X147Y121_BQ),
.O5(CLBLM_R_X93Y121_SLICE_X146Y121_DO5),
.O6(CLBLM_R_X93Y121_SLICE_X146Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0c0a0c0f0f00000)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_CLUT (
.I0(CLBLM_R_X93Y121_SLICE_X146Y121_A5Q),
.I1(CLBLM_R_X93Y121_SLICE_X147Y121_AO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X89Y122_SLICE_X140Y122_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X93Y121_SLICE_X146Y121_CO5),
.O6(CLBLM_R_X93Y121_SLICE_X146Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33ca0a0a0a0)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y121_SLICE_X146Y121_BQ),
.I2(CLBLM_R_X93Y122_SLICE_X147Y122_C5Q),
.I3(CLBLM_R_X93Y121_SLICE_X147Y121_BQ),
.I4(CLBLM_L_X92Y121_SLICE_X144Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y121_SLICE_X146Y121_BO5),
.O6(CLBLM_R_X93Y121_SLICE_X146Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X93Y121_SLICE_X146Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y121_SLICE_X146Y121_A5Q),
.I2(CLBLM_L_X92Y119_SLICE_X145Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y121_SLICE_X146Y121_AO5),
.O6(CLBLM_R_X93Y121_SLICE_X146Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X147Y121_BO5),
.Q(CLBLM_R_X93Y121_SLICE_X147Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X147Y121_CO5),
.Q(CLBLM_R_X93Y121_SLICE_X147Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X147Y121_AO5),
.Q(CLBLM_R_X93Y121_SLICE_X147Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X147Y121_BO6),
.Q(CLBLM_R_X93Y121_SLICE_X147Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y121_SLICE_X147Y121_CO6),
.Q(CLBLM_R_X93Y121_SLICE_X147Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_DLUT (
.I0(CLBLM_R_X97Y120_SLICE_X153Y120_D5Q),
.I1(CLBLM_R_X93Y121_SLICE_X147Y121_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y121_SLICE_X146Y121_CQ),
.I4(CLBLM_R_X93Y121_SLICE_X147Y121_B5Q),
.I5(CLBLM_R_X93Y121_SLICE_X147Y121_AQ),
.O5(CLBLM_R_X93Y121_SLICE_X147Y121_DO5),
.O6(CLBLM_R_X93Y121_SLICE_X147Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_CLUT (
.I0(CLBLM_R_X93Y121_SLICE_X146Y121_CQ),
.I1(1'b1),
.I2(CLBLM_L_X94Y121_SLICE_X148Y121_CQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y121_SLICE_X147Y121_CO5),
.O6(CLBLM_R_X93Y121_SLICE_X147Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X92Y121_SLICE_X144Y121_BQ),
.I2(CLBLM_R_X93Y121_SLICE_X147Y121_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y121_SLICE_X147Y121_BO5),
.O6(CLBLM_R_X93Y121_SLICE_X147Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55a88888888)
  ) CLBLM_R_X93Y121_SLICE_X147Y121_ALUT (
.I0(CLBLM_R_X93Y121_SLICE_X147Y121_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y121_SLICE_X147Y121_CQ),
.I3(CLBLM_R_X93Y121_SLICE_X147Y121_AQ),
.I4(CLBLM_R_X93Y121_SLICE_X146Y121_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y121_SLICE_X147Y121_AO5),
.O6(CLBLM_R_X93Y121_SLICE_X147Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y122_SLICE_X146Y122_AO5),
.Q(CLBLM_R_X93Y122_SLICE_X146Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y122_SLICE_X146Y122_AO6),
.Q(CLBLM_R_X93Y122_SLICE_X146Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_DO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_CO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5aa5cccca55a)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_BLUT (
.I0(CLBLM_L_X92Y123_SLICE_X145Y123_BQ),
.I1(CLBLM_R_X97Y123_SLICE_X152Y123_C5Q),
.I2(CLBLM_R_X93Y122_SLICE_X146Y122_AQ),
.I3(CLBLM_L_X92Y122_SLICE_X145Y122_B5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X92Y122_SLICE_X145Y122_AQ),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_BO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ff000000)
  ) CLBLM_R_X93Y122_SLICE_X146Y122_ALUT (
.I0(CLBLM_L_X92Y123_SLICE_X145Y123_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X93Y123_SLICE_X146Y123_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X146Y122_AO5),
.O6(CLBLM_R_X93Y122_SLICE_X146Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y122_SLICE_X147Y122_BO5),
.Q(CLBLM_R_X93Y122_SLICE_X147Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y122_SLICE_X147Y122_CO5),
.Q(CLBLM_R_X93Y122_SLICE_X147Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y122_SLICE_X147Y122_AO6),
.Q(CLBLM_R_X93Y122_SLICE_X147Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y122_SLICE_X147Y122_CO6),
.Q(CLBLM_R_X93Y122_SLICE_X147Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X93Y123_SLICE_X147Y123_C5Q),
.I2(CLBLM_R_X97Y121_SLICE_X153Y121_C5Q),
.I3(CLBLM_R_X93Y122_SLICE_X147Y122_A5Q),
.I4(CLBLM_R_X93Y122_SLICE_X147Y122_AQ),
.I5(CLBLM_R_X93Y122_SLICE_X147Y122_CQ),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_DO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y121_SLICE_X147Y121_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y122_SLICE_X147Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_CO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966c0c0c0c0)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_BLUT (
.I0(CLBLM_R_X93Y122_SLICE_X147Y122_AQ),
.I1(CLBLM_R_X93Y123_SLICE_X147Y123_C5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y122_SLICE_X147Y122_CQ),
.I4(CLBLM_R_X93Y122_SLICE_X147Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_BO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b0f0308080c000)
  ) CLBLM_R_X93Y122_SLICE_X147Y122_ALUT (
.I0(CLBLM_L_X92Y121_SLICE_X144Y121_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y122_SLICE_X147Y122_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X90Y124_SLICE_X142Y124_DO6),
.O5(CLBLM_R_X93Y122_SLICE_X147Y122_AO5),
.O6(CLBLM_R_X93Y122_SLICE_X147Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X146Y123_BO5),
.Q(CLBLM_R_X93Y123_SLICE_X146Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X146Y123_AO5),
.Q(CLBLM_R_X93Y123_SLICE_X146Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X146Y123_BO6),
.Q(CLBLM_R_X93Y123_SLICE_X146Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X147Y123_AO5),
.Q(CLBLM_R_X93Y123_SLICE_X146Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_DLUT (
.I0(CLBLM_L_X92Y123_SLICE_X144Y123_BQ),
.I1(CLBLM_R_X93Y123_SLICE_X146Y123_AQ),
.I2(CLBLM_R_X97Y123_SLICE_X153Y123_C5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X93Y123_SLICE_X146Y123_B5Q),
.I5(CLBLM_R_X93Y123_SLICE_X147Y123_BQ),
.O5(CLBLM_R_X93Y123_SLICE_X146Y123_DO5),
.O6(CLBLM_R_X93Y123_SLICE_X146Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_CLUT (
.I0(CLBLM_R_X93Y123_SLICE_X146Y123_BQ),
.I1(CLBLM_R_X93Y122_SLICE_X146Y122_A5Q),
.I2(CLBLM_R_X97Y123_SLICE_X152Y123_CQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X92Y123_SLICE_X145Y123_CQ),
.I5(CLBLM_L_X92Y123_SLICE_X145Y123_B5Q),
.O5(CLBLM_R_X93Y123_SLICE_X146Y123_CO5),
.O6(CLBLM_R_X93Y123_SLICE_X146Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_BLUT (
.I0(CLBLM_L_X92Y123_SLICE_X145Y123_CQ),
.I1(1'b1),
.I2(CLBLM_R_X93Y123_SLICE_X147Y123_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y123_SLICE_X146Y123_BO5),
.O6(CLBLM_R_X93Y123_SLICE_X146Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_R_X93Y123_SLICE_X146Y123_ALUT (
.I0(CLBLM_R_X93Y123_SLICE_X146Y123_B5Q),
.I1(CLBLM_R_X93Y123_SLICE_X146Y123_AQ),
.I2(CLBLM_R_X93Y123_SLICE_X147Y123_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y123_SLICE_X144Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y123_SLICE_X146Y123_AO5),
.O6(CLBLM_R_X93Y123_SLICE_X146Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X147Y123_BO5),
.Q(CLBLM_R_X93Y123_SLICE_X147Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X147Y123_CO5),
.Q(CLBLM_R_X93Y123_SLICE_X147Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X147Y123_BO6),
.Q(CLBLM_R_X93Y123_SLICE_X147Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y123_SLICE_X147Y123_CO6),
.Q(CLBLM_R_X93Y123_SLICE_X147Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_DLUT (
.I0(CLBLM_L_X92Y123_SLICE_X144Y123_CQ),
.I1(CLBLM_R_X93Y123_SLICE_X147Y123_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y123_SLICE_X146Y123_CQ),
.I4(CLBLM_R_X93Y123_SLICE_X147Y123_B5Q),
.I5(CLBLM_R_X97Y123_SLICE_X153Y123_CQ),
.O5(CLBLM_R_X93Y123_SLICE_X147Y123_DO5),
.O6(CLBLM_R_X93Y123_SLICE_X147Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cc00cc00)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_CLUT (
.I0(CLBLM_L_X92Y123_SLICE_X144Y123_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y122_SLICE_X147Y122_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y123_SLICE_X147Y123_CO5),
.O6(CLBLM_R_X93Y123_SLICE_X147Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c088888888)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_BLUT (
.I0(CLBLM_R_X93Y123_SLICE_X147Y123_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y123_SLICE_X144Y123_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y123_SLICE_X147Y123_BO5),
.O6(CLBLM_R_X93Y123_SLICE_X147Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f000f000)
  ) CLBLM_R_X93Y123_SLICE_X147Y123_ALUT (
.I0(CLBLM_R_X93Y123_SLICE_X147Y123_CQ),
.I1(CLBLM_R_X93Y123_SLICE_X146Y123_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y123_SLICE_X147Y123_B5Q),
.I4(CLBLM_L_X92Y123_SLICE_X144Y123_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y123_SLICE_X147Y123_AO5),
.O6(CLBLM_R_X93Y123_SLICE_X147Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X146Y124_BO5),
.Q(CLBLM_R_X93Y124_SLICE_X146Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X146Y124_CO5),
.Q(CLBLM_R_X93Y124_SLICE_X146Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X146Y124_AO6),
.Q(CLBLM_R_X93Y124_SLICE_X146Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X146Y124_CO6),
.Q(CLBLM_R_X93Y124_SLICE_X146Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_DLUT (
.I0(CLBLM_R_X93Y124_SLICE_X146Y124_C5Q),
.I1(CLBLM_R_X93Y124_SLICE_X146Y124_AQ),
.I2(CLBLM_L_X92Y122_SLICE_X144Y122_CQ),
.I3(CLBLM_R_X93Y124_SLICE_X146Y124_A5Q),
.I4(CLBLM_R_X93Y124_SLICE_X146Y124_CQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X93Y124_SLICE_X146Y124_DO5),
.O6(CLBLM_R_X93Y124_SLICE_X146Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff000000)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X93Y124_SLICE_X146Y124_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y124_SLICE_X146Y124_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y124_SLICE_X146Y124_CO5),
.O6(CLBLM_R_X93Y124_SLICE_X146Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_BLUT (
.I0(CLBLM_R_X93Y124_SLICE_X146Y124_CQ),
.I1(CLBLM_R_X93Y124_SLICE_X146Y124_A5Q),
.I2(CLBLM_R_X93Y124_SLICE_X146Y124_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y124_SLICE_X146Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y124_SLICE_X146Y124_BO5),
.O6(CLBLM_R_X93Y124_SLICE_X146Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacafa0a00000000)
  ) CLBLM_R_X93Y124_SLICE_X146Y124_ALUT (
.I0(CLBLM_R_X95Y125_SLICE_X150Y125_DO6),
.I1(CLBLM_R_X93Y126_SLICE_X146Y126_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y124_SLICE_X146Y124_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X93Y124_SLICE_X146Y124_AO5),
.O6(CLBLM_R_X93Y124_SLICE_X146Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X147Y124_AO5),
.Q(CLBLM_R_X93Y124_SLICE_X147Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X147Y124_BO5),
.Q(CLBLM_R_X93Y124_SLICE_X147Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X147Y124_CO5),
.Q(CLBLM_R_X93Y124_SLICE_X147Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X147Y124_AO6),
.Q(CLBLM_R_X93Y124_SLICE_X147Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X147Y124_BO6),
.Q(CLBLM_R_X93Y124_SLICE_X147Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y124_SLICE_X147Y124_CO6),
.Q(CLBLM_R_X93Y124_SLICE_X147Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_DLUT (
.I0(CLBLM_R_X93Y124_SLICE_X147Y124_C5Q),
.I1(CLBLM_R_X93Y124_SLICE_X147Y124_CQ),
.I2(CLBLM_R_X93Y124_SLICE_X147Y124_BQ),
.I3(1'b1),
.I4(CLBLM_R_X95Y124_SLICE_X150Y124_CQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X93Y124_SLICE_X147Y124_DO5),
.O6(CLBLM_R_X93Y124_SLICE_X147Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y124_SLICE_X147Y124_BQ),
.I4(CLBLM_R_X93Y124_SLICE_X147Y124_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y124_SLICE_X147Y124_CO5),
.O6(CLBLM_R_X93Y124_SLICE_X147Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888c0c0c0c0)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_BLUT (
.I0(CLBLM_R_X95Y124_SLICE_X150Y124_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X94Y124_SLICE_X148Y124_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y124_SLICE_X147Y124_BO5),
.O6(CLBLM_R_X93Y124_SLICE_X147Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h444444440cc0c00c)
  ) CLBLM_R_X93Y124_SLICE_X147Y124_ALUT (
.I0(CLBLM_R_X93Y120_SLICE_X146Y120_CO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y120_SLICE_X146Y120_A5Q),
.I3(CLBLM_L_X94Y124_SLICE_X148Y124_C5Q),
.I4(CLBLM_R_X93Y124_SLICE_X147Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y124_SLICE_X147Y124_AO5),
.O6(CLBLM_R_X93Y124_SLICE_X147Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y125_SLICE_X146Y125_BO5),
.Q(CLBLM_R_X93Y125_SLICE_X146Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y125_SLICE_X146Y125_CO5),
.Q(CLBLM_R_X93Y125_SLICE_X146Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y125_SLICE_X146Y125_AO6),
.Q(CLBLM_R_X93Y125_SLICE_X146Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y125_SLICE_X146Y125_CO6),
.Q(CLBLM_R_X93Y125_SLICE_X146Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_DLUT (
.I0(CLBLM_R_X93Y125_SLICE_X146Y125_C5Q),
.I1(CLBLM_R_X93Y125_SLICE_X146Y125_CQ),
.I2(CLBLM_R_X93Y125_SLICE_X146Y125_AQ),
.I3(CLBLM_R_X93Y125_SLICE_X146Y125_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X90Y124_SLICE_X143Y124_C5Q),
.O5(CLBLM_R_X93Y125_SLICE_X146Y125_DO5),
.O6(CLBLM_R_X93Y125_SLICE_X146Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff000000)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X93Y125_SLICE_X146Y125_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y125_SLICE_X146Y125_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y125_SLICE_X146Y125_CO5),
.O6(CLBLM_R_X93Y125_SLICE_X146Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_BLUT (
.I0(CLBLM_R_X93Y125_SLICE_X146Y125_CQ),
.I1(CLBLM_R_X93Y125_SLICE_X146Y125_A5Q),
.I2(CLBLM_R_X93Y125_SLICE_X146Y125_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X93Y125_SLICE_X146Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y125_SLICE_X146Y125_BO5),
.O6(CLBLM_R_X93Y125_SLICE_X146Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8fc3000000000)
  ) CLBLM_R_X93Y125_SLICE_X146Y125_ALUT (
.I0(CLBLM_R_X93Y126_SLICE_X146Y126_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X94Y125_SLICE_X148Y125_DO6),
.I3(CLBLM_R_X93Y125_SLICE_X146Y125_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X93Y125_SLICE_X146Y125_AO5),
.O6(CLBLM_R_X93Y125_SLICE_X146Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y125_SLICE_X147Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y125_SLICE_X147Y125_AO5),
.Q(CLBLM_R_X93Y125_SLICE_X147Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y125_SLICE_X147Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y125_SLICE_X147Y125_AO6),
.Q(CLBLM_R_X93Y125_SLICE_X147Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y125_SLICE_X147Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y125_SLICE_X147Y125_DO5),
.O6(CLBLM_R_X93Y125_SLICE_X147Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y125_SLICE_X147Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y125_SLICE_X147Y125_CO5),
.O6(CLBLM_R_X93Y125_SLICE_X147Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y125_SLICE_X147Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y125_SLICE_X147Y125_BO5),
.O6(CLBLM_R_X93Y125_SLICE_X147Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0000cc84848484)
  ) CLBLM_R_X93Y125_SLICE_X147Y125_ALUT (
.I0(CLBLM_R_X93Y125_SLICE_X146Y125_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y125_SLICE_X147Y125_AQ),
.I3(CLBLM_L_X92Y125_SLICE_X145Y125_A5Q),
.I4(CLBLM_R_X93Y128_SLICE_X147Y128_DQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y125_SLICE_X147Y125_AO5),
.O6(CLBLM_R_X93Y125_SLICE_X147Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X146Y126_AO5),
.Q(CLBLM_R_X93Y126_SLICE_X146Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X146Y126_CO5),
.Q(CLBLM_R_X93Y126_SLICE_X146Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X146Y126_AO6),
.Q(CLBLM_R_X93Y126_SLICE_X146Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X146Y126_BO5),
.Q(CLBLM_R_X93Y126_SLICE_X146Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X146Y126_CO6),
.Q(CLBLM_R_X93Y126_SLICE_X146Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_DLUT (
.I0(CLBLM_R_X93Y126_SLICE_X146Y126_C5Q),
.I1(CLBLM_R_X93Y126_SLICE_X146Y126_CQ),
.I2(CLBLM_R_X93Y126_SLICE_X146Y126_BQ),
.I3(CLBLM_R_X93Y129_SLICE_X146Y129_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X92Y126_SLICE_X145Y126_C5Q),
.O5(CLBLM_R_X93Y126_SLICE_X146Y126_DO5),
.O6(CLBLM_R_X93Y126_SLICE_X146Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y126_SLICE_X146Y126_CQ),
.I2(CLBLM_R_X93Y129_SLICE_X146Y129_CQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y126_SLICE_X146Y126_CO5),
.O6(CLBLM_R_X93Y126_SLICE_X146Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_BLUT (
.I0(CLBLM_R_X93Y126_SLICE_X146Y126_CQ),
.I1(CLBLM_R_X93Y126_SLICE_X146Y126_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y129_SLICE_X146Y129_CQ),
.I4(CLBLM_R_X93Y126_SLICE_X146Y126_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y126_SLICE_X146Y126_BO5),
.O6(CLBLM_R_X93Y126_SLICE_X146Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X93Y126_SLICE_X146Y126_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y127_SLICE_X146Y127_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y126_SLICE_X146Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y126_SLICE_X146Y126_AO5),
.O6(CLBLM_R_X93Y126_SLICE_X146Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X147Y126_BO5),
.Q(CLBLM_R_X93Y126_SLICE_X147Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X147Y126_CO5),
.Q(CLBLM_R_X93Y126_SLICE_X147Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X147Y126_AO6),
.Q(CLBLM_R_X93Y126_SLICE_X147Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y126_SLICE_X147Y126_CO6),
.Q(CLBLM_R_X93Y126_SLICE_X147Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_DLUT (
.I0(CLBLM_R_X93Y126_SLICE_X147Y126_C5Q),
.I1(CLBLM_R_X93Y126_SLICE_X147Y126_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y126_SLICE_X147Y126_A5Q),
.I4(CLBLM_R_X93Y126_SLICE_X147Y126_AQ),
.I5(CLBLM_L_X90Y125_SLICE_X143Y125_BQ),
.O5(CLBLM_R_X93Y126_SLICE_X147Y126_DO5),
.O6(CLBLM_R_X93Y126_SLICE_X147Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y126_SLICE_X147Y126_CQ),
.I2(CLBLM_R_X93Y126_SLICE_X147Y126_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y126_SLICE_X147Y126_CO5),
.O6(CLBLM_R_X93Y126_SLICE_X147Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996cccc0000)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_BLUT (
.I0(CLBLM_R_X93Y126_SLICE_X147Y126_CQ),
.I1(CLBLM_R_X93Y126_SLICE_X147Y126_C5Q),
.I2(CLBLM_R_X93Y126_SLICE_X147Y126_AQ),
.I3(CLBLM_R_X93Y126_SLICE_X147Y126_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X93Y126_SLICE_X147Y126_BO5),
.O6(CLBLM_R_X93Y126_SLICE_X147Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacafa0a00000000)
  ) CLBLM_R_X93Y126_SLICE_X147Y126_ALUT (
.I0(CLBLM_R_X95Y129_SLICE_X150Y129_DO6),
.I1(CLBLM_L_X94Y125_SLICE_X148Y125_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X93Y126_SLICE_X147Y126_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X93Y126_SLICE_X147Y126_AO5),
.O6(CLBLM_R_X93Y126_SLICE_X147Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y127_SLICE_X146Y127_AO5),
.Q(CLBLM_R_X93Y127_SLICE_X146Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y127_SLICE_X146Y127_AO6),
.Q(CLBLM_R_X93Y127_SLICE_X146Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y127_SLICE_X146Y127_BO6),
.Q(CLBLM_R_X93Y127_SLICE_X146Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y127_SLICE_X146Y127_CO6),
.Q(CLBLM_R_X93Y127_SLICE_X146Y127_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y127_SLICE_X146Y127_DO5),
.O6(CLBLM_R_X93Y127_SLICE_X146Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d80000ff000000)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X93Y129_SLICE_X146Y129_B5Q),
.I2(CLBLM_L_X92Y126_SLICE_X145Y126_AO6),
.I3(CLBLM_R_X95Y128_SLICE_X151Y128_AO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X93Y127_SLICE_X146Y127_CO5),
.O6(CLBLM_R_X93Y127_SLICE_X146Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b07030c0804000)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y127_SLICE_X145Y127_AO6),
.I4(CLBLM_R_X93Y130_SLICE_X146Y130_AQ),
.I5(CLBLM_R_X95Y128_SLICE_X150Y128_CO6),
.O5(CLBLM_R_X93Y127_SLICE_X146Y127_BO5),
.O6(CLBLM_R_X93Y127_SLICE_X146Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X93Y127_SLICE_X146Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y127_SLICE_X146Y127_A5Q),
.I2(CLBLM_R_X93Y130_SLICE_X146Y130_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y127_SLICE_X146Y127_AO5),
.O6(CLBLM_R_X93Y127_SLICE_X146Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y127_SLICE_X147Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y127_SLICE_X147Y127_DO5),
.O6(CLBLM_R_X93Y127_SLICE_X147Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y127_SLICE_X147Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y127_SLICE_X147Y127_CO5),
.O6(CLBLM_R_X93Y127_SLICE_X147Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y127_SLICE_X147Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y127_SLICE_X147Y127_BO5),
.O6(CLBLM_R_X93Y127_SLICE_X147Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y127_SLICE_X147Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y127_SLICE_X147Y127_AO5),
.O6(CLBLM_R_X93Y127_SLICE_X147Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X146Y128_BO5),
.Q(CLBLM_R_X93Y128_SLICE_X146Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X146Y128_CO5),
.Q(CLBLM_R_X93Y128_SLICE_X146Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X146Y128_AO6),
.Q(CLBLM_R_X93Y128_SLICE_X146Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X146Y128_CO6),
.Q(CLBLM_R_X93Y128_SLICE_X146Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000069966996)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_DLUT (
.I0(CLBLM_R_X93Y128_SLICE_X146Y128_C5Q),
.I1(CLBLM_R_X93Y128_SLICE_X146Y128_CQ),
.I2(CLBLM_R_X93Y128_SLICE_X146Y128_AQ),
.I3(CLBLM_R_X93Y128_SLICE_X146Y128_A5Q),
.I4(CLBLM_L_X90Y125_SLICE_X143Y125_DQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X93Y128_SLICE_X146Y128_DO5),
.O6(CLBLM_R_X93Y128_SLICE_X146Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X93Y128_SLICE_X146Y128_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y128_SLICE_X146Y128_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y128_SLICE_X146Y128_CO5),
.O6(CLBLM_R_X93Y128_SLICE_X146Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_BLUT (
.I0(CLBLM_R_X93Y128_SLICE_X146Y128_CQ),
.I1(CLBLM_R_X93Y128_SLICE_X146Y128_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y128_SLICE_X146Y128_AQ),
.I4(CLBLM_R_X93Y128_SLICE_X146Y128_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y128_SLICE_X146Y128_BO5),
.O6(CLBLM_R_X93Y128_SLICE_X146Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e02020e020e020)
  ) CLBLM_R_X93Y128_SLICE_X146Y128_ALUT (
.I0(CLBLM_L_X94Y128_SLICE_X149Y128_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y128_SLICE_X146Y128_BO6),
.I4(CLBLM_R_X93Y127_SLICE_X146Y127_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X93Y128_SLICE_X146Y128_AO5),
.O6(CLBLM_R_X93Y128_SLICE_X146Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X147Y128_AO5),
.Q(CLBLM_R_X93Y128_SLICE_X147Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X147Y128_BO5),
.Q(CLBLM_R_X93Y128_SLICE_X147Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X147Y128_AO6),
.Q(CLBLM_R_X93Y128_SLICE_X147Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X147Y128_BO6),
.Q(CLBLM_R_X93Y128_SLICE_X147Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X147Y128_CO6),
.Q(CLBLM_R_X93Y128_SLICE_X147Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y128_SLICE_X147Y128_DO6),
.Q(CLBLM_R_X93Y128_SLICE_X147Y128_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cccc00cc0000cc)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y120_SLICE_X146Y120_A5Q),
.I4(CLBLM_R_X93Y128_SLICE_X147Y128_CQ),
.I5(CLBLM_R_X93Y128_SLICE_X146Y128_A5Q),
.O5(CLBLM_R_X93Y128_SLICE_X147Y128_DO5),
.O6(CLBLM_R_X93Y128_SLICE_X147Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c00c0cc0c00c0c)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X92Y127_SLICE_X145Y127_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y131_SLICE_X147Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y128_SLICE_X147Y128_CO5),
.O6(CLBLM_R_X93Y128_SLICE_X147Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha050a050c0c03030)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_BLUT (
.I0(CLBLM_L_X92Y126_SLICE_X144Y126_AQ),
.I1(CLBLM_R_X93Y128_SLICE_X147Y128_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y128_SLICE_X147Y128_AQ),
.I4(CLBLM_R_X93Y126_SLICE_X146Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y128_SLICE_X147Y128_BO5),
.O6(CLBLM_R_X93Y128_SLICE_X147Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9090909050a0a050)
  ) CLBLM_R_X93Y128_SLICE_X147Y128_ALUT (
.I0(CLBLM_R_X93Y120_SLICE_X146Y120_A5Q),
.I1(CLBLM_R_X93Y126_SLICE_X147Y126_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y128_SLICE_X145Y128_A5Q),
.I4(CLBLM_R_X93Y129_SLICE_X147Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y128_SLICE_X147Y128_AO5),
.O6(CLBLM_R_X93Y128_SLICE_X147Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X146Y129_AO5),
.Q(CLBLM_R_X93Y129_SLICE_X146Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X146Y129_BO5),
.Q(CLBLM_R_X93Y129_SLICE_X146Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X146Y129_AO6),
.Q(CLBLM_R_X93Y129_SLICE_X146Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X146Y129_BO6),
.Q(CLBLM_R_X93Y129_SLICE_X146Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X146Y129_CO6),
.Q(CLBLM_R_X93Y129_SLICE_X146Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X146Y129_DO5),
.O6(CLBLM_R_X93Y129_SLICE_X146Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha088aa88a0880088)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y130_SLICE_X151Y130_DO6),
.I2(CLBLM_R_X93Y129_SLICE_X146Y129_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X93Y126_SLICE_X146Y126_BO6),
.O5(CLBLM_R_X93Y129_SLICE_X146Y129_CO5),
.O6(CLBLM_R_X93Y129_SLICE_X146Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_BLUT (
.I0(CLBLM_R_X93Y129_SLICE_X146Y129_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X94Y125_SLICE_X148Y125_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X146Y129_BO5),
.O6(CLBLM_R_X93Y129_SLICE_X146Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_R_X93Y129_SLICE_X146Y129_ALUT (
.I0(CLBLM_R_X93Y129_SLICE_X146Y129_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y129_SLICE_X146Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X146Y129_AO5),
.O6(CLBLM_R_X93Y129_SLICE_X146Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X147Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X147Y129_AO5),
.Q(CLBLM_R_X93Y129_SLICE_X147Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y129_SLICE_X147Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y129_SLICE_X147Y129_AO6),
.Q(CLBLM_R_X93Y129_SLICE_X147Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y129_SLICE_X147Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X147Y129_DO5),
.O6(CLBLM_R_X93Y129_SLICE_X147Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y129_SLICE_X147Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X147Y129_CO5),
.O6(CLBLM_R_X93Y129_SLICE_X147Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y129_SLICE_X147Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X147Y129_BO5),
.O6(CLBLM_R_X93Y129_SLICE_X147Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc003300a500a500)
  ) CLBLM_R_X93Y129_SLICE_X147Y129_ALUT (
.I0(CLBLM_R_X93Y128_SLICE_X147Y128_A5Q),
.I1(CLBLM_R_X93Y128_SLICE_X147Y128_B5Q),
.I2(CLBLM_R_X93Y131_SLICE_X146Y131_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X92Y129_SLICE_X145Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y129_SLICE_X147Y129_AO5),
.O6(CLBLM_R_X93Y129_SLICE_X147Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X146Y130_AO5),
.Q(CLBLM_R_X93Y130_SLICE_X146Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X146Y130_BO5),
.Q(CLBLM_R_X93Y130_SLICE_X146Y130_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X146Y130_AO6),
.Q(CLBLM_R_X93Y130_SLICE_X146Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X146Y130_BO6),
.Q(CLBLM_R_X93Y130_SLICE_X146Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y130_SLICE_X146Y130_DO5),
.O6(CLBLM_R_X93Y130_SLICE_X146Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y130_SLICE_X146Y130_CO5),
.O6(CLBLM_R_X93Y130_SLICE_X146Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cc00cc00)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_BLUT (
.I0(CLBLM_R_X93Y130_SLICE_X146Y130_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X93Y129_SLICE_X146Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y130_SLICE_X146Y130_BO5),
.O6(CLBLM_R_X93Y130_SLICE_X146Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X93Y130_SLICE_X146Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y130_SLICE_X146Y130_A5Q),
.I2(CLBLM_R_X93Y132_SLICE_X146Y132_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y130_SLICE_X146Y130_AO5),
.O6(CLBLM_R_X93Y130_SLICE_X146Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X147Y130_BO5),
.Q(CLBLM_R_X93Y130_SLICE_X147Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X147Y130_CO5),
.Q(CLBLM_R_X93Y130_SLICE_X147Y130_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X147Y130_AO6),
.Q(CLBLM_R_X93Y130_SLICE_X147Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y130_SLICE_X147Y130_CO6),
.Q(CLBLM_R_X93Y130_SLICE_X147Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_DLUT (
.I0(CLBLM_R_X93Y130_SLICE_X147Y130_C5Q),
.I1(CLBLM_R_X93Y130_SLICE_X147Y130_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y130_SLICE_X147Y130_A5Q),
.I4(CLBLM_R_X93Y130_SLICE_X147Y130_AQ),
.I5(CLBLM_L_X92Y131_SLICE_X144Y131_C5Q),
.O5(CLBLM_R_X93Y130_SLICE_X147Y130_DO5),
.O6(CLBLM_R_X93Y130_SLICE_X147Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y130_SLICE_X147Y130_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y130_SLICE_X147Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y130_SLICE_X147Y130_CO5),
.O6(CLBLM_R_X93Y130_SLICE_X147Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acccc0000)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_BLUT (
.I0(CLBLM_R_X93Y130_SLICE_X147Y130_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X93Y130_SLICE_X147Y130_AQ),
.I3(CLBLM_R_X93Y130_SLICE_X147Y130_A5Q),
.I4(CLBLM_R_X93Y130_SLICE_X147Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y130_SLICE_X147Y130_BO5),
.O6(CLBLM_R_X93Y130_SLICE_X147Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000cc00aa00cc00)
  ) CLBLM_R_X93Y130_SLICE_X147Y130_ALUT (
.I0(CLBLM_R_X93Y130_SLICE_X147Y130_BO6),
.I1(CLBLM_R_X95Y130_SLICE_X150Y130_DO6),
.I2(CLBLM_R_X93Y130_SLICE_X146Y130_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X93Y130_SLICE_X147Y130_AO5),
.O6(CLBLM_R_X93Y130_SLICE_X147Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X146Y131_BO5),
.Q(CLBLM_R_X93Y131_SLICE_X146Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X146Y131_CO5),
.Q(CLBLM_R_X93Y131_SLICE_X146Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X146Y131_AO6),
.Q(CLBLM_R_X93Y131_SLICE_X146Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X146Y131_CO6),
.Q(CLBLM_R_X93Y131_SLICE_X146Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f9f9f606090906)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_DLUT (
.I0(CLBLM_R_X93Y131_SLICE_X146Y131_C5Q),
.I1(CLBLM_R_X93Y131_SLICE_X146Y131_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y131_SLICE_X146Y131_A5Q),
.I4(CLBLM_R_X93Y131_SLICE_X146Y131_CQ),
.I5(CLBLM_L_X90Y128_SLICE_X143Y128_D5Q),
.O5(CLBLM_R_X93Y131_SLICE_X146Y131_DO5),
.O6(CLBLM_R_X93Y131_SLICE_X146Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X93Y131_SLICE_X146Y131_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y131_SLICE_X146Y131_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y131_SLICE_X146Y131_CO5),
.O6(CLBLM_R_X93Y131_SLICE_X146Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_BLUT (
.I0(CLBLM_R_X93Y131_SLICE_X146Y131_CQ),
.I1(CLBLM_R_X93Y131_SLICE_X146Y131_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y131_SLICE_X146Y131_A5Q),
.I4(CLBLM_R_X93Y131_SLICE_X146Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y131_SLICE_X146Y131_BO5),
.O6(CLBLM_R_X93Y131_SLICE_X146Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c0a0a03000a0a0)
  ) CLBLM_R_X93Y131_SLICE_X146Y131_ALUT (
.I0(CLBLM_R_X97Y131_SLICE_X152Y131_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y131_SLICE_X146Y131_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X93Y130_SLICE_X146Y130_B5Q),
.O5(CLBLM_R_X93Y131_SLICE_X146Y131_AO5),
.O6(CLBLM_R_X93Y131_SLICE_X146Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X147Y131_AO5),
.Q(CLBLM_R_X93Y131_SLICE_X147Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X147Y131_BO5),
.Q(CLBLM_R_X93Y131_SLICE_X147Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X147Y131_AO6),
.Q(CLBLM_R_X93Y131_SLICE_X147Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y131_SLICE_X147Y131_BO6),
.Q(CLBLM_R_X93Y131_SLICE_X147Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y131_SLICE_X147Y131_DO5),
.O6(CLBLM_R_X93Y131_SLICE_X147Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y131_SLICE_X147Y131_CO5),
.O6(CLBLM_R_X93Y131_SLICE_X147Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_BLUT (
.I0(CLBLM_R_X93Y130_SLICE_X147Y130_A5Q),
.I1(CLBLM_R_X93Y131_SLICE_X147Y131_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X92Y132_SLICE_X145Y132_A5Q),
.I4(CLBLM_R_X93Y131_SLICE_X147Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X93Y131_SLICE_X147Y131_BO5),
.O6(CLBLM_R_X93Y131_SLICE_X147Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc330000a5a50000)
  ) CLBLM_R_X93Y131_SLICE_X147Y131_ALUT (
.I0(CLBLM_R_X93Y133_SLICE_X146Y133_A5Q),
.I1(CLBLM_L_X92Y131_SLICE_X145Y131_A5Q),
.I2(CLBLM_R_X93Y131_SLICE_X147Y131_AQ),
.I3(CLBLM_R_X93Y129_SLICE_X147Y129_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X93Y131_SLICE_X147Y131_AO5),
.O6(CLBLM_R_X93Y131_SLICE_X147Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y132_SLICE_X146Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y132_SLICE_X146Y132_AO5),
.Q(CLBLM_R_X93Y132_SLICE_X146Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y132_SLICE_X146Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y132_SLICE_X146Y132_AO6),
.Q(CLBLM_R_X93Y132_SLICE_X146Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X146Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X146Y132_DO5),
.O6(CLBLM_R_X93Y132_SLICE_X146Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X146Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X146Y132_CO5),
.O6(CLBLM_R_X93Y132_SLICE_X146Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X146Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X146Y132_BO5),
.O6(CLBLM_R_X93Y132_SLICE_X146Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X93Y132_SLICE_X146Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X93Y132_SLICE_X146Y132_A5Q),
.I2(CLBLM_R_X93Y130_SLICE_X146Y130_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X146Y132_AO5),
.O6(CLBLM_R_X93Y132_SLICE_X146Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X147Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X147Y132_DO5),
.O6(CLBLM_R_X93Y132_SLICE_X147Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X147Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X147Y132_CO5),
.O6(CLBLM_R_X93Y132_SLICE_X147Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X147Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X147Y132_BO5),
.O6(CLBLM_R_X93Y132_SLICE_X147Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y132_SLICE_X147Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y132_SLICE_X147Y132_AO5),
.O6(CLBLM_R_X93Y132_SLICE_X147Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y133_SLICE_X146Y133_BO5),
.Q(CLBLM_R_X93Y133_SLICE_X146Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y133_SLICE_X146Y133_CO5),
.Q(CLBLM_R_X93Y133_SLICE_X146Y133_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y133_SLICE_X146Y133_AO6),
.Q(CLBLM_R_X93Y133_SLICE_X146Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X93Y133_SLICE_X146Y133_CO6),
.Q(CLBLM_R_X93Y133_SLICE_X146Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_DLUT (
.I0(CLBLM_R_X93Y133_SLICE_X146Y133_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X93Y133_SLICE_X146Y133_AQ),
.I3(CLBLM_R_X93Y133_SLICE_X146Y133_A5Q),
.I4(CLBLM_R_X93Y133_SLICE_X146Y133_CQ),
.I5(CLBLM_L_X92Y131_SLICE_X144Y131_B5Q),
.O5(CLBLM_R_X93Y133_SLICE_X146Y133_DO5),
.O6(CLBLM_R_X93Y133_SLICE_X146Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X93Y133_SLICE_X146Y133_AQ),
.I3(1'b1),
.I4(CLBLM_R_X93Y133_SLICE_X146Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X93Y133_SLICE_X146Y133_CO5),
.O6(CLBLM_R_X93Y133_SLICE_X146Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996cccc0000)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_BLUT (
.I0(CLBLM_R_X93Y133_SLICE_X146Y133_CQ),
.I1(CLBLM_R_X93Y133_SLICE_X146Y133_C5Q),
.I2(CLBLM_R_X93Y133_SLICE_X146Y133_AQ),
.I3(CLBLM_R_X93Y133_SLICE_X146Y133_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X93Y133_SLICE_X146Y133_BO5),
.O6(CLBLM_R_X93Y133_SLICE_X146Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7b30000c4800000)
  ) CLBLM_R_X93Y133_SLICE_X146Y133_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X93Y132_SLICE_X146Y132_A5Q),
.I3(CLBLM_R_X93Y133_SLICE_X146Y133_BO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_L_X94Y132_SLICE_X149Y132_AO6),
.O5(CLBLM_R_X93Y133_SLICE_X146Y133_AO5),
.O6(CLBLM_R_X93Y133_SLICE_X146Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y133_SLICE_X147Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y133_SLICE_X147Y133_DO5),
.O6(CLBLM_R_X93Y133_SLICE_X147Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y133_SLICE_X147Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y133_SLICE_X147Y133_CO5),
.O6(CLBLM_R_X93Y133_SLICE_X147Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y133_SLICE_X147Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y133_SLICE_X147Y133_BO5),
.O6(CLBLM_R_X93Y133_SLICE_X147Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X93Y133_SLICE_X147Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X93Y133_SLICE_X147Y133_AO5),
.O6(CLBLM_R_X93Y133_SLICE_X147Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X150Y111_AO5),
.Q(CLBLM_R_X95Y111_SLICE_X150Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X150Y111_BO5),
.Q(CLBLM_R_X95Y111_SLICE_X150Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X150Y111_CO5),
.Q(CLBLM_R_X95Y111_SLICE_X150Y111_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X150Y111_AO6),
.Q(CLBLM_R_X95Y111_SLICE_X150Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X150Y111_BO6),
.Q(CLBLM_R_X95Y111_SLICE_X150Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X150Y111_CO6),
.Q(CLBLM_R_X95Y111_SLICE_X150Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_DLUT (
.I0(CLBLM_R_X95Y111_SLICE_X150Y111_BQ),
.I1(CLBLM_R_X95Y111_SLICE_X150Y111_CQ),
.I2(CLBLM_R_X95Y111_SLICE_X150Y111_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X94Y112_SLICE_X149Y112_BQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y111_SLICE_X150Y111_DO5),
.O6(CLBLM_R_X95Y111_SLICE_X150Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_CLUT (
.I0(CLBLM_R_X95Y111_SLICE_X150Y111_BQ),
.I1(CLBLM_R_X95Y111_SLICE_X150Y111_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y111_SLICE_X150Y111_CO5),
.O6(CLBLM_R_X95Y111_SLICE_X150Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cc00cc00)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_L_X94Y111_SLICE_X149Y111_B5Q),
.I4(CLBLM_L_X94Y112_SLICE_X149Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y111_SLICE_X150Y111_BO5),
.O6(CLBLM_R_X95Y111_SLICE_X150Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500f0000f00)
  ) CLBLM_R_X95Y111_SLICE_X150Y111_ALUT (
.I0(CLBLM_R_X95Y112_SLICE_X150Y112_DO6),
.I1(1'b1),
.I2(CLBLM_R_X97Y111_SLICE_X152Y111_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y111_SLICE_X150Y111_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y111_SLICE_X150Y111_AO5),
.O6(CLBLM_R_X95Y111_SLICE_X150Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X151Y111_AO5),
.Q(CLBLM_R_X95Y111_SLICE_X151Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X151Y111_BO5),
.Q(CLBLM_R_X95Y111_SLICE_X151Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X151Y111_AO6),
.Q(CLBLM_R_X95Y111_SLICE_X151Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y111_SLICE_X151Y111_BO6),
.Q(CLBLM_R_X95Y111_SLICE_X151Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y111_SLICE_X151Y111_DO5),
.O6(CLBLM_R_X95Y111_SLICE_X151Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y113_SLICE_X150Y113_BQ),
.I2(CLBLM_R_X95Y111_SLICE_X151Y111_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X95Y111_SLICE_X151Y111_B5Q),
.I5(CLBLM_R_X95Y111_SLICE_X151Y111_AQ),
.O5(CLBLM_R_X95Y111_SLICE_X151Y111_CO5),
.O6(CLBLM_R_X95Y111_SLICE_X151Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y111_SLICE_X151Y111_BQ),
.I2(CLBLM_R_X95Y111_SLICE_X151Y111_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y111_SLICE_X151Y111_BO5),
.O6(CLBLM_R_X95Y111_SLICE_X151Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X95Y111_SLICE_X151Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y113_SLICE_X150Y113_BQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y113_SLICE_X151Y113_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y111_SLICE_X151Y111_AO5),
.O6(CLBLM_R_X95Y111_SLICE_X151Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y112_SLICE_X150Y112_AO5),
.Q(CLBLM_R_X95Y112_SLICE_X150Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y112_SLICE_X150Y112_BO5),
.Q(CLBLM_R_X95Y112_SLICE_X150Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y112_SLICE_X150Y112_AO6),
.Q(CLBLM_R_X95Y112_SLICE_X150Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y112_SLICE_X150Y112_BO6),
.Q(CLBLM_R_X95Y112_SLICE_X150Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5c0f005c5cfff0)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_DLUT (
.I0(CLBLM_R_X97Y111_SLICE_X153Y111_AQ),
.I1(CLBLM_L_X98Y111_SLICE_X155Y111_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y112_SLICE_X146Y112_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X98Y112_SLICE_X155Y112_A5Q),
.O5(CLBLM_R_X95Y112_SLICE_X150Y112_DO5),
.O6(CLBLM_R_X95Y112_SLICE_X150Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f7f25752a7a2070)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X95Y113_SLICE_X150Y113_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y112_SLICE_X154Y112_B5Q),
.I4(CLBLM_R_X97Y112_SLICE_X152Y112_DO6),
.I5(CLBLM_R_X93Y111_SLICE_X147Y111_CO6),
.O5(CLBLM_R_X95Y112_SLICE_X150Y112_CO5),
.O6(CLBLM_R_X95Y112_SLICE_X150Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa82828282)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y111_SLICE_X147Y111_A5Q),
.I2(CLBLM_R_X95Y111_SLICE_X150Y111_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X95Y112_SLICE_X150Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X95Y112_SLICE_X150Y112_BO5),
.O6(CLBLM_R_X95Y112_SLICE_X150Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444c00cc00c)
  ) CLBLM_R_X95Y112_SLICE_X150Y112_ALUT (
.I0(CLBLM_R_X95Y113_SLICE_X150Y113_CO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y112_SLICE_X150Y112_B5Q),
.I3(CLBLM_R_X93Y111_SLICE_X147Y111_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y112_SLICE_X150Y112_AO5),
.O6(CLBLM_R_X95Y112_SLICE_X150Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y112_SLICE_X151Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y112_SLICE_X151Y112_DO5),
.O6(CLBLM_R_X95Y112_SLICE_X151Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y112_SLICE_X151Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y112_SLICE_X151Y112_CO5),
.O6(CLBLM_R_X95Y112_SLICE_X151Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y112_SLICE_X151Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y112_SLICE_X151Y112_BO5),
.O6(CLBLM_R_X95Y112_SLICE_X151Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h323ef2fe020ec2ce)
  ) CLBLM_R_X95Y112_SLICE_X151Y112_ALUT (
.I0(CLBLM_R_X93Y114_SLICE_X147Y114_CO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X97Y112_SLICE_X152Y112_A5Q),
.I4(CLBLM_R_X95Y113_SLICE_X151Y113_AQ),
.I5(CLBLM_R_X95Y111_SLICE_X151Y111_CO6),
.O5(CLBLM_R_X95Y112_SLICE_X151Y112_AO5),
.O6(CLBLM_R_X95Y112_SLICE_X151Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X150Y113_AO5),
.Q(CLBLM_R_X95Y113_SLICE_X150Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X150Y113_BO5),
.Q(CLBLM_R_X95Y113_SLICE_X150Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X150Y113_AO6),
.Q(CLBLM_R_X95Y113_SLICE_X150Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X150Y113_BO6),
.Q(CLBLM_R_X95Y113_SLICE_X150Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y113_SLICE_X150Y113_DO5),
.O6(CLBLM_R_X95Y113_SLICE_X150Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h27ff27aa27552700)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X95Y113_SLICE_X150Y113_AQ),
.I2(CLBLM_L_X98Y113_SLICE_X154Y113_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X93Y113_SLICE_X146Y113_DO6),
.I5(CLBLM_R_X97Y113_SLICE_X152Y113_BO6),
.O5(CLBLM_R_X95Y113_SLICE_X150Y113_CO5),
.O6(CLBLM_R_X95Y113_SLICE_X150Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000099990000)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_BLUT (
.I0(CLBLM_R_X95Y114_SLICE_X150Y114_A5Q),
.I1(CLBLM_L_X94Y113_SLICE_X149Y113_A5Q),
.I2(CLBLM_R_X95Y112_SLICE_X151Y112_AO6),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y113_SLICE_X150Y113_BO5),
.O6(CLBLM_R_X95Y113_SLICE_X150Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ff000000)
  ) CLBLM_R_X95Y113_SLICE_X150Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y113_SLICE_X150Y113_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X97Y111_SLICE_X153Y111_AQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y113_SLICE_X150Y113_AO5),
.O6(CLBLM_R_X95Y113_SLICE_X150Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X151Y113_AO5),
.Q(CLBLM_R_X95Y113_SLICE_X151Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X151Y113_BO5),
.Q(CLBLM_R_X95Y113_SLICE_X151Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X151Y113_AO6),
.Q(CLBLM_R_X95Y113_SLICE_X151Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y113_SLICE_X151Y113_BO6),
.Q(CLBLM_R_X95Y113_SLICE_X151Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_DLUT (
.I0(CLBLM_R_X95Y114_SLICE_X150Y114_AQ),
.I1(CLBLM_R_X95Y111_SLICE_X151Y111_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X95Y113_SLICE_X151Y113_BQ),
.I4(CLBLM_R_X95Y113_SLICE_X151Y113_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y113_SLICE_X151Y113_DO5),
.O6(CLBLM_R_X95Y113_SLICE_X151Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32ba109876fe54dc)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X94Y113_SLICE_X149Y113_CO6),
.I3(CLBLM_R_X95Y113_SLICE_X151Y113_A5Q),
.I4(CLBLM_R_X95Y113_SLICE_X151Y113_DO6),
.I5(CLBLM_R_X97Y112_SLICE_X153Y112_B5Q),
.O5(CLBLM_R_X95Y113_SLICE_X151Y113_CO5),
.O6(CLBLM_R_X95Y113_SLICE_X151Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y113_SLICE_X151Y113_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y114_SLICE_X150Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y113_SLICE_X151Y113_BO5),
.O6(CLBLM_R_X95Y113_SLICE_X151Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X95Y113_SLICE_X151Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y113_SLICE_X151Y113_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y116_SLICE_X151Y116_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y113_SLICE_X151Y113_AO5),
.O6(CLBLM_R_X95Y113_SLICE_X151Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y114_SLICE_X150Y114_AO5),
.Q(CLBLM_R_X95Y114_SLICE_X150Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y114_SLICE_X150Y114_BO5),
.Q(CLBLM_R_X95Y114_SLICE_X150Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y114_SLICE_X150Y114_CO5),
.Q(CLBLM_R_X95Y114_SLICE_X150Y114_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y114_SLICE_X150Y114_AO6),
.Q(CLBLM_R_X95Y114_SLICE_X150Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y114_SLICE_X150Y114_BO6),
.Q(CLBLM_R_X95Y114_SLICE_X150Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y114_SLICE_X150Y114_CO6),
.Q(CLBLM_R_X95Y114_SLICE_X150Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_DLUT (
.I0(CLBLM_R_X95Y114_SLICE_X150Y114_C5Q),
.I1(CLBLM_R_X95Y114_SLICE_X150Y114_CQ),
.I2(CLBLM_R_X95Y115_SLICE_X150Y115_B5Q),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X95Y114_SLICE_X150Y114_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X150Y114_DO5),
.O6(CLBLM_R_X95Y114_SLICE_X150Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y114_SLICE_X150Y114_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y115_SLICE_X150Y115_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X150Y114_CO5),
.O6(CLBLM_R_X95Y114_SLICE_X150Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X94Y114_SLICE_X149Y114_BQ),
.I3(1'b1),
.I4(CLBLM_R_X95Y114_SLICE_X150Y114_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X150Y114_BO5),
.O6(CLBLM_R_X95Y114_SLICE_X150Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88228822)
  ) CLBLM_R_X95Y114_SLICE_X150Y114_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y114_SLICE_X150Y114_B5Q),
.I2(CLBLM_R_X95Y113_SLICE_X151Y113_CO6),
.I3(CLBLM_R_X93Y120_SLICE_X147Y120_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X150Y114_AO5),
.O6(CLBLM_R_X95Y114_SLICE_X150Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y114_SLICE_X151Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X151Y114_DO5),
.O6(CLBLM_R_X95Y114_SLICE_X151Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y114_SLICE_X151Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X151Y114_CO5),
.O6(CLBLM_R_X95Y114_SLICE_X151Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y114_SLICE_X151Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X151Y114_BO5),
.O6(CLBLM_R_X95Y114_SLICE_X151Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y114_SLICE_X151Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y114_SLICE_X151Y114_AO5),
.O6(CLBLM_R_X95Y114_SLICE_X151Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y115_SLICE_X150Y115_AO5),
.Q(CLBLM_R_X95Y115_SLICE_X150Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y115_SLICE_X150Y115_BO5),
.Q(CLBLM_R_X95Y115_SLICE_X150Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y115_SLICE_X150Y115_CO5),
.Q(CLBLM_R_X95Y115_SLICE_X150Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y115_SLICE_X150Y115_AO6),
.Q(CLBLM_R_X95Y115_SLICE_X150Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y115_SLICE_X150Y115_BO6),
.Q(CLBLM_R_X95Y115_SLICE_X150Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y115_SLICE_X150Y115_CO6),
.Q(CLBLM_R_X95Y115_SLICE_X150Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_DLUT (
.I0(CLBLM_R_X95Y115_SLICE_X150Y115_C5Q),
.I1(CLBLM_R_X95Y115_SLICE_X150Y115_CQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y115_SLICE_X150Y115_BQ),
.I4(CLBLM_R_X97Y116_SLICE_X152Y116_BQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y115_SLICE_X150Y115_DO5),
.O6(CLBLM_R_X95Y115_SLICE_X150Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000cccc0000)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_CLUT (
.I0(CLBLM_R_X97Y116_SLICE_X152Y116_BQ),
.I1(CLBLM_R_X95Y115_SLICE_X150Y115_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y115_SLICE_X150Y115_CO5),
.O6(CLBLM_R_X95Y115_SLICE_X150Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a22222222)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y116_SLICE_X150Y116_BO6),
.I2(CLBLM_R_X95Y115_SLICE_X151Y115_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y115_SLICE_X150Y115_BO5),
.O6(CLBLM_R_X95Y115_SLICE_X150Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X95Y115_SLICE_X150Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y116_SLICE_X150Y116_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X93Y115_SLICE_X147Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y115_SLICE_X150Y115_AO5),
.O6(CLBLM_R_X95Y115_SLICE_X150Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y115_SLICE_X151Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y115_SLICE_X151Y115_DO5),
.O6(CLBLM_R_X95Y115_SLICE_X151Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y115_SLICE_X151Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y115_SLICE_X151Y115_CO5),
.O6(CLBLM_R_X95Y115_SLICE_X151Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y115_SLICE_X151Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y115_SLICE_X151Y115_BO5),
.O6(CLBLM_R_X95Y115_SLICE_X151Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00caf0ca0fcaffca)
  ) CLBLM_R_X95Y115_SLICE_X151Y115_ALUT (
.I0(CLBLM_R_X95Y114_SLICE_X150Y114_DO6),
.I1(CLBLM_R_X95Y115_SLICE_X150Y115_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X95Y116_SLICE_X151Y116_AQ),
.I5(CLBLM_R_X97Y115_SLICE_X153Y115_A5Q),
.O5(CLBLM_R_X95Y115_SLICE_X151Y115_AO5),
.O6(CLBLM_R_X95Y115_SLICE_X151Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y116_SLICE_X150Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y116_SLICE_X150Y116_AO5),
.Q(CLBLM_R_X95Y116_SLICE_X150Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y116_SLICE_X150Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y116_SLICE_X150Y116_AO6),
.Q(CLBLM_R_X95Y116_SLICE_X150Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y116_SLICE_X150Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y116_SLICE_X150Y116_DO5),
.O6(CLBLM_R_X95Y116_SLICE_X150Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X95Y116_SLICE_X150Y116_CLUT (
.I0(CLBLM_L_X94Y113_SLICE_X148Y113_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X95Y116_SLICE_X150Y116_AQ),
.I3(CLBLM_R_X95Y116_SLICE_X150Y116_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X95Y115_SLICE_X150Y115_A5Q),
.O5(CLBLM_R_X95Y116_SLICE_X150Y116_CO5),
.O6(CLBLM_R_X95Y116_SLICE_X150Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h232f202ce3efe0ec)
  ) CLBLM_R_X95Y116_SLICE_X150Y116_BLUT (
.I0(CLBLM_R_X95Y114_SLICE_X150Y114_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y114_SLICE_X150Y114_A5Q),
.I4(CLBLM_R_X95Y121_SLICE_X151Y121_CO6),
.I5(CLBLM_L_X94Y116_SLICE_X149Y116_B5Q),
.O5(CLBLM_R_X95Y116_SLICE_X150Y116_BO5),
.O6(CLBLM_R_X95Y116_SLICE_X150Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa0000)
  ) CLBLM_R_X95Y116_SLICE_X150Y116_ALUT (
.I0(CLBLM_R_X95Y116_SLICE_X150Y116_AQ),
.I1(1'b1),
.I2(CLBLM_L_X94Y113_SLICE_X148Y113_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y116_SLICE_X150Y116_AO5),
.O6(CLBLM_R_X95Y116_SLICE_X150Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y116_SLICE_X151Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y116_SLICE_X151Y116_AO5),
.Q(CLBLM_R_X95Y116_SLICE_X151Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y116_SLICE_X151Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y116_SLICE_X151Y116_AO6),
.Q(CLBLM_R_X95Y116_SLICE_X151Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y116_SLICE_X151Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y116_SLICE_X151Y116_DO5),
.O6(CLBLM_R_X95Y116_SLICE_X151Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y116_SLICE_X151Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y116_SLICE_X151Y116_CO5),
.O6(CLBLM_R_X95Y116_SLICE_X151Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y116_SLICE_X151Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y116_SLICE_X151Y116_BO5),
.O6(CLBLM_R_X95Y116_SLICE_X151Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X95Y116_SLICE_X151Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y116_SLICE_X151Y116_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X90Y116_SLICE_X143Y116_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y116_SLICE_X151Y116_AO5),
.O6(CLBLM_R_X95Y116_SLICE_X151Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y117_SLICE_X150Y117_AO5),
.Q(CLBLM_R_X95Y117_SLICE_X150Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y117_SLICE_X150Y117_BO5),
.Q(CLBLM_R_X95Y117_SLICE_X150Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y117_SLICE_X150Y117_CO5),
.Q(CLBLM_R_X95Y117_SLICE_X150Y117_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y117_SLICE_X150Y117_AO6),
.Q(CLBLM_R_X95Y117_SLICE_X150Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y117_SLICE_X150Y117_BO6),
.Q(CLBLM_R_X95Y117_SLICE_X150Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y117_SLICE_X150Y117_CO6),
.Q(CLBLM_R_X95Y117_SLICE_X150Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X95Y118_SLICE_X151Y118_A5Q),
.I2(CLBLM_R_X95Y117_SLICE_X150Y117_BQ),
.I3(CLBLM_R_X95Y117_SLICE_X150Y117_A5Q),
.I4(CLBLM_R_X95Y117_SLICE_X150Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X150Y117_DO5),
.O6(CLBLM_R_X95Y117_SLICE_X150Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha050a050c0c03030)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_CLUT (
.I0(CLBLM_R_X95Y118_SLICE_X150Y118_C5Q),
.I1(CLBLM_R_X95Y117_SLICE_X150Y117_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y118_SLICE_X152Y118_A5Q),
.I4(CLBLM_R_X97Y117_SLICE_X152Y117_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X150Y117_CO5),
.O6(CLBLM_R_X95Y117_SLICE_X150Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y117_SLICE_X150Y117_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y117_SLICE_X150Y117_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X150Y117_BO5),
.O6(CLBLM_R_X95Y117_SLICE_X150Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa22222222)
  ) CLBLM_R_X95Y117_SLICE_X150Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y118_SLICE_X150Y118_DO6),
.I2(1'b1),
.I3(CLBLM_L_X94Y117_SLICE_X149Y117_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X150Y117_AO5),
.O6(CLBLM_R_X95Y117_SLICE_X150Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y117_SLICE_X151Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X151Y117_DO5),
.O6(CLBLM_R_X95Y117_SLICE_X151Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y117_SLICE_X151Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X151Y117_CO5),
.O6(CLBLM_R_X95Y117_SLICE_X151Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y117_SLICE_X151Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X151Y117_BO5),
.O6(CLBLM_R_X95Y117_SLICE_X151Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y117_SLICE_X151Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y117_SLICE_X151Y117_AO5),
.O6(CLBLM_R_X95Y117_SLICE_X151Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X150Y118_AO5),
.Q(CLBLM_R_X95Y118_SLICE_X150Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X150Y118_BO5),
.Q(CLBLM_R_X95Y118_SLICE_X150Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X150Y118_CO5),
.Q(CLBLM_R_X95Y118_SLICE_X150Y118_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X150Y118_AO6),
.Q(CLBLM_R_X95Y118_SLICE_X150Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X150Y118_BO6),
.Q(CLBLM_R_X95Y118_SLICE_X150Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X150Y118_CO6),
.Q(CLBLM_R_X95Y118_SLICE_X150Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa55ffe4e4e4e4)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLL_L_X102Y121_SLICE_X161Y121_DO6),
.I2(CLBLM_R_X95Y117_SLICE_X150Y117_DO6),
.I3(CLBLM_R_X97Y119_SLICE_X152Y119_A5Q),
.I4(CLBLM_R_X95Y118_SLICE_X150Y118_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X95Y118_SLICE_X150Y118_DO5),
.O6(CLBLM_R_X95Y118_SLICE_X150Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05050c030c030)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_CLUT (
.I0(CLBLM_L_X98Y119_SLICE_X154Y119_B5Q),
.I1(CLBLM_R_X95Y118_SLICE_X150Y118_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y118_SLICE_X153Y118_AQ),
.I4(CLBLM_R_X97Y119_SLICE_X152Y119_CQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y118_SLICE_X150Y118_CO5),
.O6(CLBLM_R_X95Y118_SLICE_X150Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y121_SLICE_X156Y121_C5Q),
.I2(CLBLM_R_X95Y118_SLICE_X151Y118_A5Q),
.I3(CLBLM_L_X94Y117_SLICE_X148Y117_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y118_SLICE_X150Y118_BO5),
.O6(CLBLM_R_X95Y118_SLICE_X150Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLM_R_X95Y118_SLICE_X150Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y118_SLICE_X151Y118_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X95Y118_SLICE_X150Y118_B5Q),
.I4(CLBLM_L_X94Y118_SLICE_X148Y118_BO6),
.I5(1'b1),
.O5(CLBLM_R_X95Y118_SLICE_X150Y118_AO5),
.O6(CLBLM_R_X95Y118_SLICE_X150Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X151Y118_AO5),
.Q(CLBLM_R_X95Y118_SLICE_X151Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X151Y118_BO5),
.Q(CLBLM_R_X95Y118_SLICE_X151Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X151Y118_AO6),
.Q(CLBLM_R_X95Y118_SLICE_X151Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y118_SLICE_X151Y118_BO6),
.Q(CLBLM_R_X95Y118_SLICE_X151Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y118_SLICE_X151Y118_DO5),
.O6(CLBLM_R_X95Y118_SLICE_X151Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_CLUT (
.I0(CLBLM_R_X97Y119_SLICE_X152Y119_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X95Y118_SLICE_X151Y118_BQ),
.I3(1'b1),
.I4(CLBLM_R_X95Y118_SLICE_X151Y118_AQ),
.I5(CLBLM_R_X95Y118_SLICE_X151Y118_B5Q),
.O5(CLBLM_R_X95Y118_SLICE_X151Y118_CO5),
.O6(CLBLM_R_X95Y118_SLICE_X151Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y118_SLICE_X151Y118_BQ),
.I2(CLBLM_R_X95Y118_SLICE_X151Y118_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y118_SLICE_X151Y118_BO5),
.O6(CLBLM_R_X95Y118_SLICE_X151Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X95Y118_SLICE_X151Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y117_SLICE_X150Y117_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X97Y119_SLICE_X152Y119_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y118_SLICE_X151Y118_AO5),
.O6(CLBLM_R_X95Y118_SLICE_X151Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y119_SLICE_X150Y119_AO5),
.Q(CLBLM_R_X95Y119_SLICE_X150Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y119_SLICE_X150Y119_BO5),
.Q(CLBLM_R_X95Y119_SLICE_X150Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y119_SLICE_X150Y119_CO5),
.Q(CLBLM_R_X95Y119_SLICE_X150Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y119_SLICE_X150Y119_AO6),
.Q(CLBLM_R_X95Y119_SLICE_X150Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y119_SLICE_X150Y119_BO6),
.Q(CLBLM_R_X95Y119_SLICE_X150Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y119_SLICE_X150Y119_CO6),
.Q(CLBLM_R_X95Y119_SLICE_X150Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_DLUT (
.I0(CLBLM_R_X95Y119_SLICE_X150Y119_C5Q),
.I1(CLBLM_R_X95Y119_SLICE_X150Y119_CQ),
.I2(CLBLM_R_X95Y119_SLICE_X150Y119_BQ),
.I3(CLBLM_R_X97Y120_SLICE_X153Y120_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X150Y119_DO5),
.O6(CLBLM_R_X95Y119_SLICE_X150Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y119_SLICE_X150Y119_CQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y119_SLICE_X150Y119_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X150Y119_CO5),
.O6(CLBLM_R_X95Y119_SLICE_X150Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y120_SLICE_X153Y120_AQ),
.I2(CLBLM_R_X97Y119_SLICE_X153Y119_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X150Y119_BO5),
.O6(CLBLM_R_X95Y119_SLICE_X150Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_R_X95Y119_SLICE_X150Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y119_SLICE_X150Y119_B5Q),
.I2(CLBLM_R_X95Y118_SLICE_X150Y118_A5Q),
.I3(CLBLM_L_X94Y119_SLICE_X149Y119_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X150Y119_AO5),
.O6(CLBLM_R_X95Y119_SLICE_X150Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y119_SLICE_X151Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X151Y119_DO5),
.O6(CLBLM_R_X95Y119_SLICE_X151Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y119_SLICE_X151Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X151Y119_CO5),
.O6(CLBLM_R_X95Y119_SLICE_X151Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y119_SLICE_X151Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X151Y119_BO5),
.O6(CLBLM_R_X95Y119_SLICE_X151Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y119_SLICE_X151Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y119_SLICE_X151Y119_AO5),
.O6(CLBLM_R_X95Y119_SLICE_X151Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X150Y120_AO5),
.Q(CLBLM_R_X95Y120_SLICE_X150Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X150Y120_BO5),
.Q(CLBLM_R_X95Y120_SLICE_X150Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X150Y120_AO6),
.Q(CLBLM_R_X95Y120_SLICE_X150Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X150Y120_BO6),
.Q(CLBLM_R_X95Y120_SLICE_X150Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y120_SLICE_X150Y120_DO5),
.O6(CLBLM_R_X95Y120_SLICE_X150Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_CLUT (
.I0(CLBLM_R_X95Y122_SLICE_X150Y122_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y120_SLICE_X150Y120_BQ),
.I4(CLBLM_R_X95Y120_SLICE_X150Y120_B5Q),
.I5(CLBLM_R_X95Y122_SLICE_X150Y122_BQ),
.O5(CLBLM_R_X95Y120_SLICE_X150Y120_CO5),
.O6(CLBLM_R_X95Y120_SLICE_X150Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y120_SLICE_X150Y120_BQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y122_SLICE_X150Y122_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y120_SLICE_X150Y120_BO5),
.O6(CLBLM_R_X95Y120_SLICE_X150Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f0f00000)
  ) CLBLM_R_X95Y120_SLICE_X150Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y120_SLICE_X150Y120_A5Q),
.I2(CLBLM_R_X95Y124_SLICE_X150Y124_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y120_SLICE_X150Y120_AO5),
.O6(CLBLM_R_X95Y120_SLICE_X150Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X151Y120_AO5),
.Q(CLBLM_R_X95Y120_SLICE_X151Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X151Y120_BO5),
.Q(CLBLM_R_X95Y120_SLICE_X151Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X151Y120_AO6),
.Q(CLBLM_R_X95Y120_SLICE_X151Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y120_SLICE_X151Y120_BO6),
.Q(CLBLM_R_X95Y120_SLICE_X151Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y120_SLICE_X151Y120_DO5),
.O6(CLBLM_R_X95Y120_SLICE_X151Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y120_SLICE_X151Y120_AQ),
.I2(CLBLM_R_X95Y120_SLICE_X151Y120_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X97Y123_SLICE_X153Y123_AQ),
.I5(CLBLM_R_X95Y120_SLICE_X151Y120_B5Q),
.O5(CLBLM_R_X95Y120_SLICE_X151Y120_CO5),
.O6(CLBLM_R_X95Y120_SLICE_X151Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y120_SLICE_X151Y120_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y120_SLICE_X151Y120_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y120_SLICE_X151Y120_BO5),
.O6(CLBLM_R_X95Y120_SLICE_X151Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0c0c0c0)
  ) CLBLM_R_X95Y120_SLICE_X151Y120_ALUT (
.I0(CLBLM_R_X97Y123_SLICE_X153Y123_AQ),
.I1(CLBLM_R_X95Y121_SLICE_X151Y121_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y120_SLICE_X151Y120_AO5),
.O6(CLBLM_R_X95Y120_SLICE_X151Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y121_SLICE_X150Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y121_SLICE_X150Y121_AO5),
.Q(CLBLM_R_X95Y121_SLICE_X150Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y121_SLICE_X150Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y121_SLICE_X150Y121_AO6),
.Q(CLBLM_R_X95Y121_SLICE_X150Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ff003333f0f0)
  ) CLBLM_R_X95Y121_SLICE_X150Y121_DLUT (
.I0(CLBLM_R_X95Y124_SLICE_X150Y124_AQ),
.I1(CLBLM_L_X94Y120_SLICE_X148Y120_B5Q),
.I2(CLBLM_L_X98Y122_SLICE_X155Y122_DO6),
.I3(CLBLM_R_X95Y120_SLICE_X150Y120_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y121_SLICE_X150Y121_DO5),
.O6(CLBLM_R_X95Y121_SLICE_X150Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555f0f03333ff00)
  ) CLBLM_R_X95Y121_SLICE_X150Y121_CLUT (
.I0(CLBLM_R_X95Y120_SLICE_X150Y120_A5Q),
.I1(CLBLM_R_X95Y121_SLICE_X150Y121_AQ),
.I2(CLBLM_R_X97Y121_SLICE_X152Y121_DO6),
.I3(CLBLM_R_X97Y122_SLICE_X153Y122_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y121_SLICE_X150Y121_CO5),
.O6(CLBLM_R_X95Y121_SLICE_X150Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5140d9c87362fbea)
  ) CLBLM_R_X95Y121_SLICE_X150Y121_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X95Y121_SLICE_X151Y121_CO6),
.I3(CLBLM_R_X101Y121_SLICE_X158Y121_CO6),
.I4(CLBLM_R_X95Y120_SLICE_X150Y120_AQ),
.I5(CLBLM_R_X95Y121_SLICE_X150Y121_A5Q),
.O5(CLBLM_R_X95Y121_SLICE_X150Y121_BO5),
.O6(CLBLM_R_X95Y121_SLICE_X150Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h90909090f00000f0)
  ) CLBLM_R_X95Y121_SLICE_X150Y121_ALUT (
.I0(CLBLM_R_X97Y121_SLICE_X152Y121_B5Q),
.I1(CLBLM_L_X94Y120_SLICE_X148Y120_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y121_SLICE_X151Y121_A5Q),
.I4(CLBLM_R_X95Y121_SLICE_X150Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y121_SLICE_X150Y121_AO5),
.O6(CLBLM_R_X95Y121_SLICE_X150Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y121_SLICE_X151Y121_AO5),
.Q(CLBLM_R_X95Y121_SLICE_X151Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y121_SLICE_X151Y121_BO5),
.Q(CLBLM_R_X95Y121_SLICE_X151Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y121_SLICE_X151Y121_AO6),
.Q(CLBLM_R_X95Y121_SLICE_X151Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y121_SLICE_X151Y121_BO6),
.Q(CLBLM_R_X95Y121_SLICE_X151Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_DLUT (
.I0(CLBLM_R_X95Y121_SLICE_X151Y121_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(1'b1),
.I3(CLBLM_R_X97Y121_SLICE_X153Y121_BQ),
.I4(CLBLM_R_X95Y121_SLICE_X151Y121_B5Q),
.I5(CLBLM_R_X95Y120_SLICE_X151Y120_A5Q),
.O5(CLBLM_R_X95Y121_SLICE_X151Y121_DO5),
.O6(CLBLM_R_X95Y121_SLICE_X151Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_CLUT (
.I0(CLBLM_R_X97Y121_SLICE_X152Y121_AQ),
.I1(CLBLM_R_X97Y121_SLICE_X152Y121_BQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y121_SLICE_X151Y121_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X95Y121_SLICE_X151Y121_AQ),
.O5(CLBLM_R_X95Y121_SLICE_X151Y121_CO5),
.O6(CLBLM_R_X95Y121_SLICE_X151Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y121_SLICE_X151Y121_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X97Y121_SLICE_X153Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y121_SLICE_X151Y121_BO5),
.O6(CLBLM_R_X95Y121_SLICE_X151Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X95Y121_SLICE_X151Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y121_SLICE_X152Y121_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y121_SLICE_X151Y121_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y121_SLICE_X151Y121_AO5),
.O6(CLBLM_R_X95Y121_SLICE_X151Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y122_SLICE_X150Y122_AO5),
.Q(CLBLM_R_X95Y122_SLICE_X150Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y122_SLICE_X150Y122_BO5),
.Q(CLBLM_R_X95Y122_SLICE_X150Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y122_SLICE_X150Y122_CO5),
.Q(CLBLM_R_X95Y122_SLICE_X150Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y122_SLICE_X150Y122_AO6),
.Q(CLBLM_R_X95Y122_SLICE_X150Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y122_SLICE_X150Y122_BO6),
.Q(CLBLM_R_X95Y122_SLICE_X150Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y122_SLICE_X150Y122_CO6),
.Q(CLBLM_R_X95Y122_SLICE_X150Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_DLUT (
.I0(CLBLM_R_X95Y122_SLICE_X150Y122_C5Q),
.I1(CLBLM_R_X95Y122_SLICE_X150Y122_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X95Y122_SLICE_X150Y122_B5Q),
.I5(CLBLM_R_X95Y124_SLICE_X150Y124_BQ),
.O5(CLBLM_R_X95Y122_SLICE_X150Y122_DO5),
.O6(CLBLM_R_X95Y122_SLICE_X150Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y122_SLICE_X150Y122_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y124_SLICE_X150Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y122_SLICE_X150Y122_CO5),
.O6(CLBLM_R_X95Y122_SLICE_X150Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0f00000)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y122_SLICE_X150Y122_AQ),
.I4(CLBLM_R_X95Y122_SLICE_X150Y122_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y122_SLICE_X150Y122_BO5),
.O6(CLBLM_R_X95Y122_SLICE_X150Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f0a0a05050)
  ) CLBLM_R_X95Y122_SLICE_X150Y122_ALUT (
.I0(CLBLM_R_X95Y124_SLICE_X150Y124_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y121_SLICE_X150Y121_DO6),
.I4(CLBLM_R_X97Y123_SLICE_X152Y123_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y122_SLICE_X150Y122_AO5),
.O6(CLBLM_R_X95Y122_SLICE_X150Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y122_SLICE_X151Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y122_SLICE_X151Y122_DO5),
.O6(CLBLM_R_X95Y122_SLICE_X151Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y122_SLICE_X151Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y122_SLICE_X151Y122_CO5),
.O6(CLBLM_R_X95Y122_SLICE_X151Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y122_SLICE_X151Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y122_SLICE_X151Y122_BO5),
.O6(CLBLM_R_X95Y122_SLICE_X151Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff3a3a00f03a3a)
  ) CLBLM_R_X95Y122_SLICE_X151Y122_ALUT (
.I0(CLBLM_R_X97Y125_SLICE_X152Y125_CO6),
.I1(CLBLM_L_X94Y120_SLICE_X149Y120_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y121_SLICE_X153Y121_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X95Y120_SLICE_X151Y120_CO6),
.O5(CLBLM_R_X95Y122_SLICE_X151Y122_AO5),
.O6(CLBLM_R_X95Y122_SLICE_X151Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X150Y123_AO5),
.Q(CLBLM_R_X95Y123_SLICE_X150Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X150Y123_BO5),
.Q(CLBLM_R_X95Y123_SLICE_X150Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X150Y123_AO6),
.Q(CLBLM_R_X95Y123_SLICE_X150Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X150Y123_BO6),
.Q(CLBLM_R_X95Y123_SLICE_X150Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y123_SLICE_X150Y123_DO5),
.O6(CLBLM_R_X95Y123_SLICE_X150Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_CLUT (
.I0(CLBLM_R_X95Y123_SLICE_X150Y123_BQ),
.I1(CLBLM_R_X97Y123_SLICE_X152Y123_AQ),
.I2(1'b1),
.I3(CLBLM_R_X95Y123_SLICE_X150Y123_A5Q),
.I4(CLBLM_R_X95Y123_SLICE_X150Y123_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y123_SLICE_X150Y123_CO5),
.O6(CLBLM_R_X95Y123_SLICE_X150Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff000000)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X97Y123_SLICE_X152Y123_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y123_SLICE_X150Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y123_SLICE_X150Y123_BO5),
.O6(CLBLM_R_X95Y123_SLICE_X150Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000aa00aa00)
  ) CLBLM_R_X95Y123_SLICE_X150Y123_ALUT (
.I0(CLBLM_R_X95Y123_SLICE_X150Y123_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X97Y125_SLICE_X152Y125_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y123_SLICE_X150Y123_AO5),
.O6(CLBLM_R_X95Y123_SLICE_X150Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X151Y123_AO5),
.Q(CLBLM_R_X95Y123_SLICE_X151Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X151Y123_BO5),
.Q(CLBLM_R_X95Y123_SLICE_X151Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X151Y123_AO6),
.Q(CLBLM_R_X95Y123_SLICE_X151Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y123_SLICE_X151Y123_BO6),
.Q(CLBLM_R_X95Y123_SLICE_X151Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_DLUT (
.I0(CLBLM_R_X95Y123_SLICE_X150Y123_AQ),
.I1(1'b1),
.I2(CLBLM_R_X97Y125_SLICE_X152Y125_AQ),
.I3(CLBLM_R_X95Y123_SLICE_X151Y123_BQ),
.I4(CLBLM_R_X95Y123_SLICE_X151Y123_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y123_SLICE_X151Y123_DO5),
.O6(CLBLM_R_X95Y123_SLICE_X151Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cfc0cfc5f5f5050)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_CLUT (
.I0(CLBLM_L_X94Y122_SLICE_X149Y122_B5Q),
.I1(CLBLM_R_X95Y123_SLICE_X150Y123_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X95Y123_SLICE_X151Y123_A5Q),
.I4(CLBLM_R_X97Y125_SLICE_X153Y125_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y123_SLICE_X151Y123_CO5),
.O6(CLBLM_R_X95Y123_SLICE_X151Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_BLUT (
.I0(CLBLM_R_X95Y123_SLICE_X151Y123_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y123_SLICE_X150Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y123_SLICE_X151Y123_BO5),
.O6(CLBLM_R_X95Y123_SLICE_X151Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X95Y123_SLICE_X151Y123_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X97Y121_SLICE_X153Y121_AQ),
.I3(1'b1),
.I4(CLBLM_R_X95Y123_SLICE_X151Y123_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y123_SLICE_X151Y123_AO5),
.O6(CLBLM_R_X95Y123_SLICE_X151Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X150Y124_AO5),
.Q(CLBLM_R_X95Y124_SLICE_X150Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X150Y124_BO5),
.Q(CLBLM_R_X95Y124_SLICE_X150Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X150Y124_CO5),
.Q(CLBLM_R_X95Y124_SLICE_X150Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X150Y124_AO6),
.Q(CLBLM_R_X95Y124_SLICE_X150Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X150Y124_BO6),
.Q(CLBLM_R_X95Y124_SLICE_X150Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X150Y124_CO6),
.Q(CLBLM_R_X95Y124_SLICE_X150Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50fa50fa4444eeee)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X97Y123_SLICE_X152Y123_DO6),
.I2(CLBLM_R_X95Y122_SLICE_X150Y122_DO6),
.I3(CLBLM_R_X95Y124_SLICE_X150Y124_A5Q),
.I4(CLBLM_L_X94Y120_SLICE_X148Y120_C5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y124_SLICE_X150Y124_DO5),
.O6(CLBLM_R_X95Y124_SLICE_X150Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000f00f0000)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_CLUT (
.I0(CLBLM_L_X94Y124_SLICE_X149Y124_BO6),
.I1(1'b1),
.I2(CLBLM_L_X94Y125_SLICE_X148Y125_B5Q),
.I3(CLBLM_R_X95Y125_SLICE_X151Y125_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y124_SLICE_X150Y124_CO5),
.O6(CLBLM_R_X95Y124_SLICE_X150Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h550055003c00c300)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_BLUT (
.I0(CLBLM_R_X95Y124_SLICE_X150Y124_DO6),
.I1(CLBLM_L_X98Y125_SLICE_X154Y125_D5Q),
.I2(CLBLM_L_X94Y128_SLICE_X149Y128_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y124_SLICE_X150Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y124_SLICE_X150Y124_BO5),
.O6(CLBLM_R_X95Y124_SLICE_X150Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X95Y124_SLICE_X150Y124_ALUT (
.I0(CLBLM_L_X94Y124_SLICE_X148Y124_AQ),
.I1(CLBLM_R_X95Y124_SLICE_X150Y124_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y124_SLICE_X150Y124_AO5),
.O6(CLBLM_R_X95Y124_SLICE_X150Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X151Y124_BO5),
.Q(CLBLM_R_X95Y124_SLICE_X151Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X151Y124_CO5),
.Q(CLBLM_R_X95Y124_SLICE_X151Y124_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X151Y124_AO6),
.Q(CLBLM_R_X95Y124_SLICE_X151Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y124_SLICE_X151Y124_CO6),
.Q(CLBLM_R_X95Y124_SLICE_X151Y124_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acaca3aca3a3ac)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_DLUT (
.I0(CLBLM_L_X94Y124_SLICE_X148Y124_C5Q),
.I1(CLBLM_R_X95Y124_SLICE_X151Y124_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X95Y124_SLICE_X151Y124_A5Q),
.I4(CLBLM_R_X95Y124_SLICE_X151Y124_AQ),
.I5(CLBLM_R_X97Y124_SLICE_X152Y124_B5Q),
.O5(CLBLM_R_X95Y124_SLICE_X151Y124_DO5),
.O6(CLBLM_R_X95Y124_SLICE_X151Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X94Y125_SLICE_X149Y125_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y124_SLICE_X151Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y124_SLICE_X151Y124_CO5),
.O6(CLBLM_R_X95Y124_SLICE_X151Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55acc00cc00)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_BLUT (
.I0(CLBLM_R_X95Y124_SLICE_X151Y124_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y124_SLICE_X151Y124_AQ),
.I3(CLBLM_R_X97Y124_SLICE_X152Y124_B5Q),
.I4(CLBLM_R_X95Y124_SLICE_X151Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y124_SLICE_X151Y124_BO5),
.O6(CLBLM_R_X95Y124_SLICE_X151Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee002200e200e200)
  ) CLBLM_R_X95Y124_SLICE_X151Y124_ALUT (
.I0(CLBLL_L_X100Y124_SLICE_X156Y124_CO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X95Y124_SLICE_X151Y124_BO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y125_SLICE_X150Y125_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X95Y124_SLICE_X151Y124_AO5),
.O6(CLBLM_R_X95Y124_SLICE_X151Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y125_SLICE_X150Y125_AO5),
.Q(CLBLM_R_X95Y125_SLICE_X150Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y125_SLICE_X150Y125_CO5),
.Q(CLBLM_R_X95Y125_SLICE_X150Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y125_SLICE_X150Y125_AO6),
.Q(CLBLM_R_X95Y125_SLICE_X150Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y125_SLICE_X150Y125_BO6),
.Q(CLBLM_R_X95Y125_SLICE_X150Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_DLUT (
.I0(CLBLM_R_X95Y124_SLICE_X151Y124_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X95Y125_SLICE_X150Y125_BQ),
.I3(CLBLM_L_X94Y125_SLICE_X149Y125_CQ),
.I4(CLBLM_R_X95Y125_SLICE_X150Y125_B5Q),
.I5(CLBLM_L_X94Y124_SLICE_X148Y124_CQ),
.O5(CLBLM_R_X95Y125_SLICE_X150Y125_DO5),
.O6(CLBLM_R_X95Y125_SLICE_X150Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y125_SLICE_X150Y125_B5Q),
.I2(CLBLM_R_X95Y125_SLICE_X150Y125_BQ),
.I3(CLBLM_L_X94Y125_SLICE_X149Y125_CQ),
.I4(CLBLM_R_X95Y124_SLICE_X151Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y125_SLICE_X150Y125_CO5),
.O6(CLBLM_R_X95Y125_SLICE_X150Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd080f0a0d0805000)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X95Y125_SLICE_X150Y125_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y125_SLICE_X155Y125_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y125_SLICE_X150Y125_CO6),
.O5(CLBLM_R_X95Y125_SLICE_X150Y125_BO5),
.O6(CLBLM_R_X95Y125_SLICE_X150Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X95Y125_SLICE_X150Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y125_SLICE_X150Y125_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X94Y127_SLICE_X149Y127_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y125_SLICE_X150Y125_AO5),
.O6(CLBLM_R_X95Y125_SLICE_X150Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y125_SLICE_X151Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y125_SLICE_X151Y125_AO5),
.Q(CLBLM_R_X95Y125_SLICE_X151Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y125_SLICE_X151Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y125_SLICE_X151Y125_AO6),
.Q(CLBLM_R_X95Y125_SLICE_X151Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y125_SLICE_X151Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y125_SLICE_X151Y125_DO5),
.O6(CLBLM_R_X95Y125_SLICE_X151Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X95Y125_SLICE_X151Y125_CLUT (
.I0(CLBLM_R_X95Y126_SLICE_X150Y126_AQ),
.I1(CLBLM_R_X97Y127_SLICE_X153Y127_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y125_SLICE_X151Y125_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X95Y125_SLICE_X151Y125_AQ),
.O5(CLBLM_R_X95Y125_SLICE_X151Y125_CO5),
.O6(CLBLM_R_X95Y125_SLICE_X151Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00ffaaaacccc)
  ) CLBLM_R_X95Y125_SLICE_X151Y125_BLUT (
.I0(CLBLM_R_X95Y123_SLICE_X151Y123_DO6),
.I1(CLBLM_R_X97Y126_SLICE_X152Y126_CO6),
.I2(CLBLM_R_X95Y123_SLICE_X151Y123_AQ),
.I3(CLBLM_L_X94Y122_SLICE_X149Y122_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X95Y125_SLICE_X151Y125_BO5),
.O6(CLBLM_R_X95Y125_SLICE_X151Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f000f000)
  ) CLBLM_R_X95Y125_SLICE_X151Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y125_SLICE_X151Y125_AQ),
.I4(CLBLM_R_X95Y126_SLICE_X150Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y125_SLICE_X151Y125_AO5),
.O6(CLBLM_R_X95Y125_SLICE_X151Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y126_SLICE_X150Y126_AO5),
.Q(CLBLM_R_X95Y126_SLICE_X150Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y126_SLICE_X150Y126_BO5),
.Q(CLBLM_R_X95Y126_SLICE_X150Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y126_SLICE_X150Y126_AO6),
.Q(CLBLM_R_X95Y126_SLICE_X150Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y126_SLICE_X150Y126_BO6),
.Q(CLBLM_R_X95Y126_SLICE_X150Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y126_SLICE_X150Y126_DO5),
.O6(CLBLM_R_X95Y126_SLICE_X150Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_R_X95Y126_SLICE_X150Y126_BQ),
.I3(CLBLM_R_X95Y126_SLICE_X150Y126_A5Q),
.I4(CLBLM_R_X95Y126_SLICE_X150Y126_B5Q),
.I5(CLBLM_R_X97Y126_SLICE_X152Y126_AQ),
.O5(CLBLM_R_X95Y126_SLICE_X150Y126_CO5),
.O6(CLBLM_R_X95Y126_SLICE_X150Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_BLUT (
.I0(CLBLM_R_X95Y126_SLICE_X150Y126_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X97Y126_SLICE_X152Y126_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y126_SLICE_X150Y126_BO5),
.O6(CLBLM_R_X95Y126_SLICE_X150Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000aa00aa00)
  ) CLBLM_R_X95Y126_SLICE_X150Y126_ALUT (
.I0(CLBLM_R_X95Y126_SLICE_X150Y126_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X97Y127_SLICE_X153Y127_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y126_SLICE_X150Y126_AO5),
.O6(CLBLM_R_X95Y126_SLICE_X150Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y126_SLICE_X151Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y126_SLICE_X151Y126_AO5),
.Q(CLBLM_R_X95Y126_SLICE_X151Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y126_SLICE_X151Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y126_SLICE_X151Y126_AO6),
.Q(CLBLM_R_X95Y126_SLICE_X151Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y126_SLICE_X151Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y126_SLICE_X151Y126_DO5),
.O6(CLBLM_R_X95Y126_SLICE_X151Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y126_SLICE_X151Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y126_SLICE_X151Y126_CO5),
.O6(CLBLM_R_X95Y126_SLICE_X151Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h32023e0ef2c2fece)
  ) CLBLM_R_X95Y126_SLICE_X151Y126_BLUT (
.I0(CLBLM_R_X97Y127_SLICE_X152Y127_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X95Y126_SLICE_X150Y126_CO6),
.I4(CLBLM_L_X94Y125_SLICE_X148Y125_B5Q),
.I5(CLBLM_R_X95Y126_SLICE_X151Y126_A5Q),
.O5(CLBLM_R_X95Y126_SLICE_X151Y126_BO5),
.O6(CLBLM_R_X95Y126_SLICE_X151Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X95Y126_SLICE_X151Y126_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y126_SLICE_X151Y126_A5Q),
.I2(CLBLM_R_X95Y123_SLICE_X151Y123_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y126_SLICE_X151Y126_AO5),
.O6(CLBLM_R_X95Y126_SLICE_X151Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y128_SLICE_X150Y128_BO5),
.Q(CLBLM_R_X95Y128_SLICE_X150Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y128_SLICE_X150Y128_AO5),
.Q(CLBLM_R_X95Y128_SLICE_X150Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y128_SLICE_X150Y128_BO6),
.Q(CLBLM_R_X95Y128_SLICE_X150Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y128_SLICE_X150Y128_DO5),
.O6(CLBLM_R_X95Y128_SLICE_X150Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0069699696)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_CLUT (
.I0(CLBLM_R_X95Y130_SLICE_X150Y130_AQ),
.I1(CLBLM_R_X95Y128_SLICE_X150Y128_AQ),
.I2(CLBLM_R_X95Y130_SLICE_X150Y130_CQ),
.I3(CLBLM_R_X93Y128_SLICE_X147Y128_CQ),
.I4(CLBLM_R_X95Y128_SLICE_X150Y128_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X95Y128_SLICE_X150Y128_CO5),
.O6(CLBLM_R_X95Y128_SLICE_X150Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y130_SLICE_X150Y130_CQ),
.I3(1'b1),
.I4(CLBLM_L_X94Y127_SLICE_X149Y127_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y128_SLICE_X150Y128_BO5),
.O6(CLBLM_R_X95Y128_SLICE_X150Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696aa00aa00)
  ) CLBLM_R_X95Y128_SLICE_X150Y128_ALUT (
.I0(CLBLM_R_X95Y128_SLICE_X150Y128_B5Q),
.I1(CLBLM_R_X95Y130_SLICE_X150Y130_AQ),
.I2(CLBLM_R_X95Y128_SLICE_X150Y128_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y130_SLICE_X150Y130_CQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y128_SLICE_X150Y128_AO5),
.O6(CLBLM_R_X95Y128_SLICE_X150Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y128_SLICE_X151Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y128_SLICE_X151Y128_DO5),
.O6(CLBLM_R_X95Y128_SLICE_X151Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y128_SLICE_X151Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y128_SLICE_X151Y128_CO5),
.O6(CLBLM_R_X95Y128_SLICE_X151Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X95Y128_SLICE_X151Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y128_SLICE_X151Y128_BO5),
.O6(CLBLM_R_X95Y128_SLICE_X151Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_R_X95Y128_SLICE_X151Y128_ALUT (
.I0(CLBLM_R_X95Y129_SLICE_X151Y129_DQ),
.I1(CLBLM_R_X95Y130_SLICE_X151Y130_C5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y128_SLICE_X147Y128_BQ),
.I4(CLBLM_R_X95Y129_SLICE_X151Y129_B5Q),
.I5(CLBLM_R_X95Y129_SLICE_X151Y129_BQ),
.O5(CLBLM_R_X95Y128_SLICE_X151Y128_AO5),
.O6(CLBLM_R_X95Y128_SLICE_X151Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X150Y129_BO5),
.Q(CLBLM_R_X95Y129_SLICE_X150Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X150Y129_CO5),
.Q(CLBLM_R_X95Y129_SLICE_X150Y129_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X150Y129_AO6),
.Q(CLBLM_R_X95Y129_SLICE_X150Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X150Y129_CO6),
.Q(CLBLM_R_X95Y129_SLICE_X150Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeebebbe14414114)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X95Y129_SLICE_X150Y129_AQ),
.I2(CLBLM_R_X95Y129_SLICE_X151Y129_D5Q),
.I3(CLBLM_R_X95Y129_SLICE_X150Y129_A5Q),
.I4(CLBLM_R_X95Y129_SLICE_X150Y129_CQ),
.I5(CLBLM_R_X93Y128_SLICE_X147Y128_AQ),
.O5(CLBLM_R_X95Y129_SLICE_X150Y129_DO5),
.O6(CLBLM_R_X95Y129_SLICE_X150Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y129_SLICE_X150Y129_AQ),
.I2(CLBLM_L_X94Y129_SLICE_X148Y129_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y129_SLICE_X150Y129_CO5),
.O6(CLBLM_R_X95Y129_SLICE_X150Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696cc00cc00)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_BLUT (
.I0(CLBLM_R_X95Y129_SLICE_X150Y129_CQ),
.I1(CLBLM_R_X95Y129_SLICE_X151Y129_D5Q),
.I2(CLBLM_R_X95Y129_SLICE_X150Y129_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y129_SLICE_X150Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y129_SLICE_X150Y129_BO5),
.O6(CLBLM_R_X95Y129_SLICE_X150Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b07030c0804000)
  ) CLBLM_R_X95Y129_SLICE_X150Y129_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y129_SLICE_X150Y129_BO6),
.I4(CLBLM_R_X95Y129_SLICE_X151Y129_A5Q),
.I5(CLBLM_L_X98Y129_SLICE_X154Y129_CO6),
.O5(CLBLM_R_X95Y129_SLICE_X150Y129_AO5),
.O6(CLBLM_R_X95Y129_SLICE_X150Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X151Y129_AO5),
.Q(CLBLM_R_X95Y129_SLICE_X151Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X151Y129_CO5),
.Q(CLBLM_R_X95Y129_SLICE_X151Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X151Y129_DO5),
.Q(CLBLM_R_X95Y129_SLICE_X151Y129_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X151Y129_AO6),
.Q(CLBLM_R_X95Y129_SLICE_X151Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X151Y129_BO6),
.Q(CLBLM_R_X95Y129_SLICE_X151Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y129_SLICE_X151Y129_DO6),
.Q(CLBLM_R_X95Y129_SLICE_X151Y129_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X95Y129_SLICE_X151Y129_BQ),
.I3(CLBLM_R_X95Y129_SLICE_X150Y129_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y129_SLICE_X151Y129_DO5),
.O6(CLBLM_R_X95Y129_SLICE_X151Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55a88888888)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_CLUT (
.I0(CLBLM_R_X95Y130_SLICE_X151Y130_C5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y129_SLICE_X151Y129_BQ),
.I3(CLBLM_R_X95Y129_SLICE_X151Y129_DQ),
.I4(CLBLM_R_X95Y129_SLICE_X151Y129_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y129_SLICE_X151Y129_CO5),
.O6(CLBLM_R_X95Y129_SLICE_X151Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc088cc88c0880088)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_BLUT (
.I0(CLBLM_L_X98Y129_SLICE_X155Y129_DO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y129_SLICE_X151Y129_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y129_SLICE_X151Y129_CO6),
.O5(CLBLM_R_X95Y129_SLICE_X151Y129_BO5),
.O6(CLBLM_R_X95Y129_SLICE_X151Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c00000cccc)
  ) CLBLM_R_X95Y129_SLICE_X151Y129_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X95Y129_SLICE_X151Y129_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X95Y126_SLICE_X151Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y129_SLICE_X151Y129_AO5),
.O6(CLBLM_R_X95Y129_SLICE_X151Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X150Y130_BO5),
.Q(CLBLM_R_X95Y130_SLICE_X150Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X150Y130_CO5),
.Q(CLBLM_R_X95Y130_SLICE_X150Y130_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X150Y130_AO6),
.Q(CLBLM_R_X95Y130_SLICE_X150Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X150Y130_CO6),
.Q(CLBLM_R_X95Y130_SLICE_X150Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f06699f0f09966)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_DLUT (
.I0(CLBLM_R_X95Y130_SLICE_X150Y130_C5Q),
.I1(CLBLM_R_X95Y131_SLICE_X150Y131_CQ),
.I2(CLBLM_R_X93Y131_SLICE_X147Y131_B5Q),
.I3(CLBLM_R_X95Y130_SLICE_X150Y130_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y132_SLICE_X150Y132_BQ),
.O5(CLBLM_R_X95Y130_SLICE_X150Y130_DO5),
.O6(CLBLM_R_X95Y130_SLICE_X150Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaaa0000)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y130_SLICE_X150Y130_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y132_SLICE_X150Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y130_SLICE_X150Y130_CO5),
.O6(CLBLM_R_X95Y130_SLICE_X150Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_BLUT (
.I0(CLBLM_R_X95Y131_SLICE_X150Y131_CQ),
.I1(CLBLM_R_X95Y130_SLICE_X150Y130_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y132_SLICE_X150Y132_BQ),
.I4(CLBLM_R_X95Y130_SLICE_X150Y130_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y130_SLICE_X150Y130_BO5),
.O6(CLBLM_R_X95Y130_SLICE_X150Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he020e020e0e02020)
  ) CLBLM_R_X95Y130_SLICE_X150Y130_ALUT (
.I0(CLBLM_L_X98Y130_SLICE_X154Y130_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X94Y130_SLICE_X149Y130_A5Q),
.I4(CLBLM_R_X95Y128_SLICE_X150Y128_AO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X95Y130_SLICE_X150Y130_AO5),
.O6(CLBLM_R_X95Y130_SLICE_X150Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X151Y130_BO5),
.Q(CLBLM_R_X95Y130_SLICE_X151Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X151Y130_CO5),
.Q(CLBLM_R_X95Y130_SLICE_X151Y130_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X151Y130_AO6),
.Q(CLBLM_R_X95Y130_SLICE_X151Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y130_SLICE_X151Y130_CO6),
.Q(CLBLM_R_X95Y130_SLICE_X151Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_DLUT (
.I0(CLBLM_R_X95Y130_SLICE_X151Y130_A5Q),
.I1(CLBLM_R_X95Y130_SLICE_X151Y130_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X93Y128_SLICE_X147Y128_B5Q),
.I4(CLBLM_R_X95Y130_SLICE_X151Y130_AQ),
.I5(CLBLM_R_X95Y131_SLICE_X151Y131_D5Q),
.O5(CLBLM_R_X95Y130_SLICE_X151Y130_DO5),
.O6(CLBLM_R_X95Y130_SLICE_X151Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y129_SLICE_X151Y129_DQ),
.I2(CLBLM_R_X95Y130_SLICE_X151Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y130_SLICE_X151Y130_CO5),
.O6(CLBLM_R_X95Y130_SLICE_X151Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996ff000000)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_BLUT (
.I0(CLBLM_R_X95Y130_SLICE_X151Y130_AQ),
.I1(CLBLM_R_X95Y130_SLICE_X151Y130_A5Q),
.I2(CLBLM_R_X95Y130_SLICE_X151Y130_CQ),
.I3(CLBLM_R_X95Y131_SLICE_X151Y131_D5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X95Y130_SLICE_X151Y130_BO5),
.O6(CLBLM_R_X95Y130_SLICE_X151Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f000c0c0c0c0)
  ) CLBLM_R_X95Y130_SLICE_X151Y130_ALUT (
.I0(CLBLM_R_X95Y131_SLICE_X150Y131_B5Q),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_DO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y130_SLICE_X151Y130_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y130_SLICE_X151Y130_AO5),
.O6(CLBLM_R_X95Y130_SLICE_X151Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X150Y131_AO5),
.Q(CLBLM_R_X95Y131_SLICE_X150Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X150Y131_BO5),
.Q(CLBLM_R_X95Y131_SLICE_X150Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X150Y131_AO6),
.Q(CLBLM_R_X95Y131_SLICE_X150Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X150Y131_BO6),
.Q(CLBLM_R_X95Y131_SLICE_X150Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X150Y131_CO6),
.Q(CLBLM_R_X95Y131_SLICE_X150Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_DLUT (
.I0(CLBLM_R_X93Y129_SLICE_X147Y129_AQ),
.I1(CLBLM_R_X95Y131_SLICE_X151Y131_A5Q),
.I2(CLBLM_R_X95Y131_SLICE_X151Y131_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X95Y131_SLICE_X151Y131_DQ),
.I5(CLBLM_R_X95Y131_SLICE_X151Y131_C5Q),
.O5(CLBLM_R_X95Y131_SLICE_X150Y131_DO5),
.O6(CLBLM_R_X95Y131_SLICE_X150Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha808a808aaaa0000)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y130_SLICE_X150Y130_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X95Y132_SLICE_X151Y132_AQ),
.I4(CLBLM_R_X97Y133_SLICE_X152Y133_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y131_SLICE_X150Y131_CO5),
.O6(CLBLM_R_X95Y131_SLICE_X150Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f0f00000)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_BLUT (
.I0(CLBLM_R_X95Y131_SLICE_X150Y131_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y129_SLICE_X151Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y131_SLICE_X150Y131_BO5),
.O6(CLBLM_R_X95Y131_SLICE_X150Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_R_X95Y131_SLICE_X150Y131_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y131_SLICE_X150Y131_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y131_SLICE_X150Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y131_SLICE_X150Y131_AO5),
.O6(CLBLM_R_X95Y131_SLICE_X150Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X151Y131_BO5),
.Q(CLBLM_R_X95Y131_SLICE_X151Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X151Y131_CO5),
.Q(CLBLM_R_X95Y131_SLICE_X151Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X151Y131_DO5),
.Q(CLBLM_R_X95Y131_SLICE_X151Y131_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X151Y131_AO6),
.Q(CLBLM_R_X95Y131_SLICE_X151Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X151Y131_CO6),
.Q(CLBLM_R_X95Y131_SLICE_X151Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y131_SLICE_X151Y131_DO6),
.Q(CLBLM_R_X95Y131_SLICE_X151Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y130_SLICE_X151Y130_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y131_SLICE_X151Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y131_SLICE_X151Y131_DO5),
.O6(CLBLM_R_X95Y131_SLICE_X151Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X95Y131_SLICE_X151Y131_DQ),
.I3(CLBLM_R_X97Y131_SLICE_X153Y131_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y131_SLICE_X151Y131_CO5),
.O6(CLBLM_R_X95Y131_SLICE_X151Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966f0f00000)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_BLUT (
.I0(CLBLM_R_X95Y131_SLICE_X151Y131_AQ),
.I1(CLBLM_R_X95Y131_SLICE_X151Y131_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y131_SLICE_X151Y131_DQ),
.I4(CLBLM_R_X95Y131_SLICE_X151Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y131_SLICE_X151Y131_BO5),
.O6(CLBLM_R_X95Y131_SLICE_X151Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f000c0c0c0c0)
  ) CLBLM_R_X95Y131_SLICE_X151Y131_ALUT (
.I0(CLBLM_R_X95Y131_SLICE_X150Y131_BQ),
.I1(CLBLM_R_X97Y131_SLICE_X153Y131_DO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y131_SLICE_X151Y131_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X95Y131_SLICE_X151Y131_AO5),
.O6(CLBLM_R_X95Y131_SLICE_X151Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X150Y132_BO5),
.Q(CLBLM_R_X95Y132_SLICE_X150Y132_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X150Y132_CO5),
.Q(CLBLM_R_X95Y132_SLICE_X150Y132_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X150Y132_AO5),
.Q(CLBLM_R_X95Y132_SLICE_X150Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X150Y132_BO6),
.Q(CLBLM_R_X95Y132_SLICE_X150Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X150Y132_CO6),
.Q(CLBLM_R_X95Y132_SLICE_X150Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_DLUT (
.I0(CLBLM_R_X93Y131_SLICE_X147Y131_BQ),
.I1(CLBLM_R_X95Y132_SLICE_X150Y132_CQ),
.I2(CLBLM_R_X95Y132_SLICE_X150Y132_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X95Y132_SLICE_X150Y132_B5Q),
.I5(CLBLM_R_X95Y132_SLICE_X151Y132_BQ),
.O5(CLBLM_R_X95Y132_SLICE_X150Y132_DO5),
.O6(CLBLM_R_X95Y132_SLICE_X150Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y132_SLICE_X152Y132_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X95Y132_SLICE_X151Y132_BQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y132_SLICE_X150Y132_CO5),
.O6(CLBLM_R_X95Y132_SLICE_X150Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0a0a0a0a0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_BLUT (
.I0(CLBLM_R_X95Y132_SLICE_X150Y132_CQ),
.I1(CLBLM_R_X95Y131_SLICE_X150Y131_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y132_SLICE_X150Y132_BO5),
.O6(CLBLM_R_X95Y132_SLICE_X150Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966c0c0c0c0)
  ) CLBLM_R_X95Y132_SLICE_X150Y132_ALUT (
.I0(CLBLM_R_X95Y132_SLICE_X150Y132_CQ),
.I1(CLBLM_R_X95Y132_SLICE_X150Y132_B5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y132_SLICE_X151Y132_BQ),
.I4(CLBLM_R_X95Y132_SLICE_X150Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X95Y132_SLICE_X150Y132_AO5),
.O6(CLBLM_R_X95Y132_SLICE_X150Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X151Y132_AO5),
.Q(CLBLM_R_X95Y132_SLICE_X151Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X151Y132_DO5),
.Q(CLBLM_R_X95Y132_SLICE_X151Y132_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X151Y132_AO6),
.Q(CLBLM_R_X95Y132_SLICE_X151Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X151Y132_BO6),
.Q(CLBLM_R_X95Y132_SLICE_X151Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X95Y132_SLICE_X151Y132_CO6),
.Q(CLBLM_R_X95Y132_SLICE_X151Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caa00aa00)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_DLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y132_SLICE_X151Y132_CQ),
.I2(CLBLM_R_X97Y132_SLICE_X152Y132_DQ),
.I3(CLBLM_R_X95Y132_SLICE_X150Y132_C5Q),
.I4(CLBLM_R_X95Y132_SLICE_X151Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X95Y132_SLICE_X151Y132_DO5),
.O6(CLBLM_R_X95Y132_SLICE_X151Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0d08070205000)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y134_SLICE_X154Y134_DO6),
.I4(CLBLM_R_X95Y132_SLICE_X151Y132_DO6),
.I5(CLBLM_R_X97Y132_SLICE_X152Y132_AQ),
.O5(CLBLM_R_X95Y132_SLICE_X151Y132_CO5),
.O6(CLBLM_R_X95Y132_SLICE_X151Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaa000030aa0000)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_BLUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X95Y132_SLICE_X150Y132_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X95Y132_SLICE_X151Y132_A5Q),
.O5(CLBLM_R_X95Y132_SLICE_X151Y132_BO5),
.O6(CLBLM_R_X95Y132_SLICE_X151Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X95Y132_SLICE_X151Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X95Y132_SLICE_X151Y132_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y132_SLICE_X152Y132_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X95Y132_SLICE_X151Y132_AO5),
.O6(CLBLM_R_X95Y132_SLICE_X151Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y111_SLICE_X152Y111_AO5),
.Q(CLBLM_R_X97Y111_SLICE_X152Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y111_SLICE_X152Y111_BO5),
.Q(CLBLM_R_X97Y111_SLICE_X152Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y111_SLICE_X152Y111_AO6),
.Q(CLBLM_R_X97Y111_SLICE_X152Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y111_SLICE_X152Y111_BO6),
.Q(CLBLM_R_X97Y111_SLICE_X152Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_DLUT (
.I0(CLBLM_R_X97Y111_SLICE_X152Y111_BQ),
.I1(CLBLM_R_X97Y111_SLICE_X152Y111_AQ),
.I2(CLBLM_L_X98Y111_SLICE_X155Y111_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X97Y111_SLICE_X152Y111_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y111_SLICE_X152Y111_DO5),
.O6(CLBLM_R_X97Y111_SLICE_X152Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7750225077fa22fa)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X97Y111_SLICE_X153Y111_A5Q),
.I2(CLBLM_R_X95Y111_SLICE_X150Y111_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X97Y111_SLICE_X152Y111_DO6),
.I5(CLBLM_L_X98Y111_SLICE_X155Y111_A5Q),
.O5(CLBLM_R_X97Y111_SLICE_X152Y111_CO5),
.O6(CLBLM_R_X97Y111_SLICE_X152Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y111_SLICE_X152Y111_BQ),
.I2(CLBLM_R_X97Y111_SLICE_X152Y111_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y111_SLICE_X152Y111_BO5),
.O6(CLBLM_R_X97Y111_SLICE_X152Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLM_R_X97Y111_SLICE_X152Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y112_SLICE_X152Y112_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X95Y111_SLICE_X150Y111_B5Q),
.I4(CLBLM_R_X97Y111_SLICE_X152Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X97Y111_SLICE_X152Y111_AO5),
.O6(CLBLM_R_X97Y111_SLICE_X152Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y111_SLICE_X153Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y111_SLICE_X153Y111_AO5),
.Q(CLBLM_R_X97Y111_SLICE_X153Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y111_SLICE_X153Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y111_SLICE_X153Y111_AO6),
.Q(CLBLM_R_X97Y111_SLICE_X153Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y111_SLICE_X153Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y111_SLICE_X153Y111_DO5),
.O6(CLBLM_R_X97Y111_SLICE_X153Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y111_SLICE_X153Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y111_SLICE_X153Y111_CO5),
.O6(CLBLM_R_X97Y111_SLICE_X153Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0faa0faa33ff3300)
  ) CLBLM_R_X97Y111_SLICE_X153Y111_BLUT (
.I0(CLBLM_L_X98Y111_SLICE_X154Y111_CO6),
.I1(CLBLL_L_X100Y111_SLICE_X157Y111_B5Q),
.I2(CLBLM_R_X97Y112_SLICE_X153Y112_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X94Y111_SLICE_X149Y111_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y111_SLICE_X153Y111_BO5),
.O6(CLBLM_R_X97Y111_SLICE_X153Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y111_SLICE_X153Y111_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y111_SLICE_X153Y111_A5Q),
.I2(CLBLM_R_X97Y112_SLICE_X153Y112_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y111_SLICE_X153Y111_AO5),
.O6(CLBLM_R_X97Y111_SLICE_X153Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X152Y112_AO5),
.Q(CLBLM_R_X97Y112_SLICE_X152Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X152Y112_BO5),
.Q(CLBLM_R_X97Y112_SLICE_X152Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X152Y112_CO5),
.Q(CLBLM_R_X97Y112_SLICE_X152Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X152Y112_AO6),
.Q(CLBLM_R_X97Y112_SLICE_X152Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X152Y112_BO6),
.Q(CLBLM_R_X97Y112_SLICE_X152Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X152Y112_CO6),
.Q(CLBLM_R_X97Y112_SLICE_X152Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_DLUT (
.I0(CLBLM_R_X97Y112_SLICE_X152Y112_C5Q),
.I1(CLBLM_R_X97Y112_SLICE_X152Y112_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X97Y112_SLICE_X152Y112_B5Q),
.I5(CLBLM_R_X95Y112_SLICE_X150Y112_BQ),
.O5(CLBLM_R_X97Y112_SLICE_X152Y112_DO5),
.O6(CLBLM_R_X97Y112_SLICE_X152Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y112_SLICE_X152Y112_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y112_SLICE_X150Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y112_SLICE_X152Y112_CO5),
.O6(CLBLM_R_X97Y112_SLICE_X152Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X95Y112_SLICE_X150Y112_AQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y112_SLICE_X152Y112_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y112_SLICE_X152Y112_BO5),
.O6(CLBLM_R_X97Y112_SLICE_X152Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaa00aa00a)
  ) CLBLM_R_X97Y112_SLICE_X152Y112_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y112_SLICE_X153Y112_B5Q),
.I3(CLBLM_R_X95Y111_SLICE_X151Y111_B5Q),
.I4(CLBLM_R_X97Y111_SLICE_X153Y111_BO6),
.I5(1'b1),
.O5(CLBLM_R_X97Y112_SLICE_X152Y112_AO5),
.O6(CLBLM_R_X97Y112_SLICE_X152Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X153Y112_AO5),
.Q(CLBLM_R_X97Y112_SLICE_X153Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X153Y112_BO5),
.Q(CLBLM_R_X97Y112_SLICE_X153Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X153Y112_AO6),
.Q(CLBLM_R_X97Y112_SLICE_X153Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y112_SLICE_X153Y112_BO6),
.Q(CLBLM_R_X97Y112_SLICE_X153Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y112_SLICE_X153Y112_DO5),
.O6(CLBLM_R_X97Y112_SLICE_X153Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff00f05c5c5c5c)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_CLUT (
.I0(CLBLL_L_X100Y111_SLICE_X157Y111_C5Q),
.I1(CLBLM_R_X95Y111_SLICE_X151Y111_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y112_SLICE_X153Y112_A5Q),
.I4(CLBLM_L_X98Y110_SLICE_X154Y110_BO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y112_SLICE_X153Y112_CO5),
.O6(CLBLM_R_X97Y112_SLICE_X153Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa88228822)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y111_SLICE_X151Y111_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X97Y115_SLICE_X153Y115_A5Q),
.I4(CLBLM_R_X97Y112_SLICE_X153Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X97Y112_SLICE_X153Y112_BO5),
.O6(CLBLM_R_X97Y112_SLICE_X153Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X97Y112_SLICE_X153Y112_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y112_SLICE_X153Y112_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y115_SLICE_X154Y115_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y112_SLICE_X153Y112_AO5),
.O6(CLBLM_R_X97Y112_SLICE_X153Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y113_SLICE_X152Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y113_SLICE_X152Y113_AO5),
.Q(CLBLM_R_X97Y113_SLICE_X152Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y113_SLICE_X152Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y113_SLICE_X152Y113_AO6),
.Q(CLBLM_R_X97Y113_SLICE_X152Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y113_SLICE_X152Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X152Y113_DO5),
.O6(CLBLM_R_X97Y113_SLICE_X152Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y113_SLICE_X152Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X152Y113_CO5),
.O6(CLBLM_R_X97Y113_SLICE_X152Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y113_SLICE_X152Y113_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y112_SLICE_X152Y112_BQ),
.I2(CLBLM_R_X97Y113_SLICE_X152Y113_AQ),
.I3(1'b1),
.I4(CLBLM_R_X95Y112_SLICE_X150Y112_AQ),
.I5(CLBLM_R_X97Y113_SLICE_X152Y113_A5Q),
.O5(CLBLM_R_X97Y113_SLICE_X152Y113_BO5),
.O6(CLBLM_R_X97Y113_SLICE_X152Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X97Y113_SLICE_X152Y113_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y113_SLICE_X152Y113_AQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y112_SLICE_X152Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X152Y113_AO5),
.O6(CLBLM_R_X97Y113_SLICE_X152Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y113_SLICE_X153Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X153Y113_DO5),
.O6(CLBLM_R_X97Y113_SLICE_X153Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y113_SLICE_X153Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X153Y113_CO5),
.O6(CLBLM_R_X97Y113_SLICE_X153Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y113_SLICE_X153Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X153Y113_BO5),
.O6(CLBLM_R_X97Y113_SLICE_X153Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y113_SLICE_X153Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y113_SLICE_X153Y113_AO5),
.O6(CLBLM_R_X97Y113_SLICE_X153Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y115_SLICE_X152Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y115_SLICE_X152Y115_AO5),
.Q(CLBLM_R_X97Y115_SLICE_X152Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y115_SLICE_X152Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y115_SLICE_X152Y115_AO6),
.Q(CLBLM_R_X97Y115_SLICE_X152Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y115_SLICE_X152Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y115_SLICE_X152Y115_DO5),
.O6(CLBLM_R_X97Y115_SLICE_X152Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y115_SLICE_X152Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y115_SLICE_X152Y115_CO5),
.O6(CLBLM_R_X97Y115_SLICE_X152Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y115_SLICE_X152Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y115_SLICE_X152Y115_BO5),
.O6(CLBLM_R_X97Y115_SLICE_X152Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88228822)
  ) CLBLM_R_X97Y115_SLICE_X152Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y115_SLICE_X148Y115_A5Q),
.I2(CLBLM_L_X98Y116_SLICE_X154Y116_AO6),
.I3(CLBLM_L_X98Y114_SLICE_X154Y114_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y115_SLICE_X152Y115_AO5),
.O6(CLBLM_R_X97Y115_SLICE_X152Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y115_SLICE_X153Y115_AO5),
.Q(CLBLM_R_X97Y115_SLICE_X153Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y115_SLICE_X153Y115_BO5),
.Q(CLBLM_R_X97Y115_SLICE_X153Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y115_SLICE_X153Y115_AO6),
.Q(CLBLM_R_X97Y115_SLICE_X153Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y115_SLICE_X153Y115_BO6),
.Q(CLBLM_R_X97Y115_SLICE_X153Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y116_SLICE_X153Y116_AQ),
.I2(CLBLM_R_X97Y115_SLICE_X153Y115_BQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y115_SLICE_X153Y115_B5Q),
.I5(CLBLM_R_X97Y116_SLICE_X153Y116_BQ),
.O5(CLBLM_R_X97Y115_SLICE_X153Y115_DO5),
.O6(CLBLM_R_X97Y115_SLICE_X153Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30fa300a3ffa3f0a)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_CLUT (
.I0(CLBLM_R_X97Y116_SLICE_X153Y116_DO6),
.I1(CLBLM_L_X98Y115_SLICE_X155Y115_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y115_SLICE_X153Y115_DO6),
.I5(CLBLL_L_X100Y115_SLICE_X156Y115_C5Q),
.O5(CLBLM_R_X97Y115_SLICE_X153Y115_CO5),
.O6(CLBLM_R_X97Y115_SLICE_X153Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y115_SLICE_X153Y115_BQ),
.I2(1'b1),
.I3(CLBLM_R_X97Y116_SLICE_X153Y116_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y115_SLICE_X153Y115_BO5),
.O6(CLBLM_R_X97Y115_SLICE_X153Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_R_X97Y115_SLICE_X153Y115_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y116_SLICE_X152Y116_A5Q),
.I2(CLBLM_R_X95Y115_SLICE_X150Y115_C5Q),
.I3(CLBLM_L_X98Y113_SLICE_X154Y113_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y115_SLICE_X153Y115_AO5),
.O6(CLBLM_R_X97Y115_SLICE_X153Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X152Y116_AO5),
.Q(CLBLM_R_X97Y116_SLICE_X152Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X152Y116_BO5),
.Q(CLBLM_R_X97Y116_SLICE_X152Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X152Y116_AO6),
.Q(CLBLM_R_X97Y116_SLICE_X152Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X152Y116_BO6),
.Q(CLBLM_R_X97Y116_SLICE_X152Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X152Y116_DO5),
.O6(CLBLM_R_X97Y116_SLICE_X152Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h333300fff0f0aaaa)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_CLUT (
.I0(CLBLM_R_X93Y120_SLICE_X147Y120_DO6),
.I1(CLBLM_R_X95Y116_SLICE_X151Y116_A5Q),
.I2(CLBLM_R_X97Y116_SLICE_X153Y116_DO6),
.I3(CLBLM_R_X97Y116_SLICE_X152Y116_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X97Y116_SLICE_X152Y116_CO5),
.O6(CLBLM_R_X97Y116_SLICE_X152Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y116_SLICE_X153Y116_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X95Y115_SLICE_X150Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X152Y116_BO5),
.O6(CLBLM_R_X97Y116_SLICE_X152Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000099990000)
  ) CLBLM_R_X97Y116_SLICE_X152Y116_ALUT (
.I0(CLBLM_R_X97Y116_SLICE_X152Y116_B5Q),
.I1(CLBLM_L_X90Y116_SLICE_X143Y116_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y115_SLICE_X154Y115_CO6),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X152Y116_AO5),
.O6(CLBLM_R_X97Y116_SLICE_X152Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X153Y116_AO5),
.Q(CLBLM_R_X97Y116_SLICE_X153Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X153Y116_BO5),
.Q(CLBLM_R_X97Y116_SLICE_X153Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X153Y116_CO5),
.Q(CLBLM_R_X97Y116_SLICE_X153Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X153Y116_AO6),
.Q(CLBLM_R_X97Y116_SLICE_X153Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X153Y116_BO6),
.Q(CLBLM_R_X97Y116_SLICE_X153Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y116_SLICE_X153Y116_CO6),
.Q(CLBLM_R_X97Y116_SLICE_X153Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_DLUT (
.I0(CLBLM_R_X97Y116_SLICE_X153Y116_C5Q),
.I1(CLBLM_R_X97Y116_SLICE_X153Y116_CQ),
.I2(CLBLM_R_X97Y116_SLICE_X152Y116_B5Q),
.I3(CLBLM_R_X97Y116_SLICE_X153Y116_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X153Y116_DO5),
.O6(CLBLM_R_X97Y116_SLICE_X153Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y116_SLICE_X153Y116_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y116_SLICE_X153Y116_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X153Y116_CO5),
.O6(CLBLM_R_X97Y116_SLICE_X153Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y116_SLICE_X155Y116_B5Q),
.I3(CLBLM_R_X97Y116_SLICE_X153Y116_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X153Y116_BO5),
.O6(CLBLM_R_X97Y116_SLICE_X153Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa0a0a0a0a)
  ) CLBLM_R_X97Y116_SLICE_X153Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y116_SLICE_X152Y116_CO6),
.I3(CLBLM_R_X97Y115_SLICE_X153Y115_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y116_SLICE_X153Y116_AO5),
.O6(CLBLM_R_X97Y116_SLICE_X153Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X152Y117_AO5),
.Q(CLBLM_R_X97Y117_SLICE_X152Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X153Y117_DO6),
.Q(CLBLM_R_X97Y117_SLICE_X152Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X152Y117_AO6),
.Q(CLBLM_R_X97Y117_SLICE_X152Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X152Y117_BO6),
.Q(CLBLM_R_X97Y117_SLICE_X152Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_DLUT (
.I0(CLBLM_R_X97Y117_SLICE_X153Y117_CQ),
.I1(CLBLM_R_X93Y117_SLICE_X146Y117_AQ),
.I2(CLBLM_R_X97Y117_SLICE_X152Y117_AQ),
.I3(CLBLM_R_X97Y117_SLICE_X152Y117_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y117_SLICE_X152Y117_DO5),
.O6(CLBLM_R_X97Y117_SLICE_X152Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff550033f033f0)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_CLUT (
.I0(CLBLM_R_X97Y117_SLICE_X153Y117_AQ),
.I1(CLBLM_R_X97Y117_SLICE_X152Y117_BQ),
.I2(CLBLM_R_X89Y115_SLICE_X141Y115_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y117_SLICE_X152Y117_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y117_SLICE_X152Y117_CO5),
.O6(CLBLM_R_X97Y117_SLICE_X152Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0aa0a0a0a00a0a)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y118_SLICE_X157Y118_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X95Y117_SLICE_X150Y117_C5Q),
.I5(CLBLM_R_X97Y117_SLICE_X152Y117_A5Q),
.O5(CLBLM_R_X97Y117_SLICE_X152Y117_BO5),
.O6(CLBLM_R_X97Y117_SLICE_X152Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y117_SLICE_X152Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y117_SLICE_X153Y117_CQ),
.I2(CLBLM_R_X97Y117_SLICE_X152Y117_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y117_SLICE_X152Y117_AO5),
.O6(CLBLM_R_X97Y117_SLICE_X152Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X153Y117_AO5),
.Q(CLBLM_R_X97Y117_SLICE_X153Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X153Y117_CO5),
.Q(CLBLM_R_X97Y117_SLICE_X153Y117_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X153Y117_AO6),
.Q(CLBLM_R_X97Y117_SLICE_X153Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X153Y117_BO6),
.Q(CLBLM_R_X97Y117_SLICE_X153Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y117_SLICE_X153Y117_CO6),
.Q(CLBLM_R_X97Y117_SLICE_X153Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a066999966)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_DLUT (
.I0(CLBLM_R_X97Y117_SLICE_X153Y117_C5Q),
.I1(CLBLM_R_X97Y117_SLICE_X153Y117_BQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y117_SLICE_X152Y117_B5Q),
.I4(CLBLM_R_X97Y118_SLICE_X153Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y117_SLICE_X153Y117_DO5),
.O6(CLBLM_R_X97Y117_SLICE_X153Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0f00000)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X93Y117_SLICE_X146Y117_AQ),
.I4(CLBLM_R_X97Y118_SLICE_X153Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y117_SLICE_X153Y117_CO5),
.O6(CLBLM_R_X97Y117_SLICE_X153Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa288802a220800)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y117_SLICE_X153Y117_DO5),
.I4(CLBLM_L_X90Y116_SLICE_X142Y116_DO6),
.I5(CLBLM_R_X97Y117_SLICE_X153Y117_A5Q),
.O5(CLBLM_R_X97Y117_SLICE_X153Y117_BO5),
.O6(CLBLM_R_X97Y117_SLICE_X153Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y117_SLICE_X153Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y117_SLICE_X153Y117_A5Q),
.I2(CLBLM_R_X97Y119_SLICE_X153Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y117_SLICE_X153Y117_AO5),
.O6(CLBLM_R_X97Y117_SLICE_X153Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X152Y118_BO5),
.Q(CLBLM_R_X97Y118_SLICE_X152Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X152Y118_CO5),
.Q(CLBLM_R_X97Y118_SLICE_X152Y118_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X152Y118_AO6),
.Q(CLBLM_R_X97Y118_SLICE_X152Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X152Y118_CO6),
.Q(CLBLM_R_X97Y118_SLICE_X152Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006969ff009696)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_DLUT (
.I0(CLBLM_R_X97Y118_SLICE_X152Y118_A5Q),
.I1(CLBLM_R_X97Y118_SLICE_X152Y118_AQ),
.I2(CLBLM_R_X97Y118_SLICE_X153Y118_B5Q),
.I3(CLBLL_L_X100Y118_SLICE_X157Y118_CQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X97Y118_SLICE_X152Y118_CQ),
.O5(CLBLM_R_X97Y118_SLICE_X152Y118_DO5),
.O6(CLBLM_R_X97Y118_SLICE_X152Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y118_SLICE_X152Y118_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y118_SLICE_X153Y118_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y118_SLICE_X152Y118_CO5),
.O6(CLBLM_R_X97Y118_SLICE_X152Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c88888888)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y118_SLICE_X153Y118_B5Q),
.I2(CLBLM_R_X97Y118_SLICE_X152Y118_AQ),
.I3(CLBLM_R_X97Y118_SLICE_X152Y118_CQ),
.I4(CLBLM_R_X97Y118_SLICE_X152Y118_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y118_SLICE_X152Y118_BO5),
.O6(CLBLM_R_X97Y118_SLICE_X152Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa882200a0a0a0a0)
  ) CLBLM_R_X97Y118_SLICE_X152Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_L_X90Y117_SLICE_X142Y117_DO6),
.I3(CLBLM_R_X97Y118_SLICE_X152Y118_BO6),
.I4(CLBLM_R_X97Y119_SLICE_X153Y119_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y118_SLICE_X152Y118_AO5),
.O6(CLBLM_R_X97Y118_SLICE_X152Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X153Y118_BO5),
.Q(CLBLM_R_X97Y118_SLICE_X153Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X153Y118_CO5),
.Q(CLBLM_R_X97Y118_SLICE_X153Y118_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X153Y118_AO5),
.Q(CLBLM_R_X97Y118_SLICE_X153Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X153Y118_BO6),
.Q(CLBLM_R_X97Y118_SLICE_X153Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y118_SLICE_X153Y118_CO6),
.Q(CLBLM_R_X97Y118_SLICE_X153Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14eb41eb41be14)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X97Y118_SLICE_X153Y118_CQ),
.I2(CLBLM_R_X97Y119_SLICE_X153Y119_BQ),
.I3(CLBLL_L_X100Y118_SLICE_X157Y118_B5Q),
.I4(CLBLM_R_X97Y118_SLICE_X153Y118_AQ),
.I5(CLBLM_R_X97Y118_SLICE_X152Y118_C5Q),
.O5(CLBLM_R_X97Y118_SLICE_X153Y118_DO5),
.O6(CLBLM_R_X97Y118_SLICE_X153Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0f00000)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y119_SLICE_X153Y119_BQ),
.I4(CLBLM_L_X98Y120_SLICE_X154Y120_CQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y118_SLICE_X153Y118_CO5),
.O6(CLBLM_R_X97Y118_SLICE_X153Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y118_SLICE_X152Y118_CQ),
.I2(CLBLM_R_X97Y117_SLICE_X153Y117_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y118_SLICE_X153Y118_BO5),
.O6(CLBLM_R_X97Y118_SLICE_X153Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996ff000000)
  ) CLBLM_R_X97Y118_SLICE_X153Y118_ALUT (
.I0(CLBLM_R_X97Y118_SLICE_X153Y118_CQ),
.I1(CLBLM_R_X97Y119_SLICE_X153Y119_BQ),
.I2(CLBLM_R_X97Y118_SLICE_X153Y118_AQ),
.I3(CLBLM_R_X97Y118_SLICE_X152Y118_C5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y118_SLICE_X153Y118_AO5),
.O6(CLBLM_R_X97Y118_SLICE_X153Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X152Y119_AO5),
.Q(CLBLM_R_X97Y119_SLICE_X152Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X152Y119_BO5),
.Q(CLBLM_R_X97Y119_SLICE_X152Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X152Y119_AO6),
.Q(CLBLM_R_X97Y119_SLICE_X152Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X152Y119_BO6),
.Q(CLBLM_R_X97Y119_SLICE_X152Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X152Y119_CO6),
.Q(CLBLM_R_X97Y119_SLICE_X152Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e4e55004e4effaa)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X95Y118_SLICE_X151Y118_CO6),
.I2(CLBLM_R_X97Y119_SLICE_X152Y119_AQ),
.I3(CLBLM_L_X98Y119_SLICE_X155Y119_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X95Y118_SLICE_X150Y118_A5Q),
.O5(CLBLM_R_X97Y119_SLICE_X152Y119_DO5),
.O6(CLBLM_R_X97Y119_SLICE_X152Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6090609060906090)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_CLUT (
.I0(CLBLL_L_X100Y119_SLICE_X156Y119_AQ),
.I1(CLBLL_L_X100Y118_SLICE_X157Y118_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y120_SLICE_X152Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y119_SLICE_X152Y119_CO5),
.O6(CLBLM_R_X97Y119_SLICE_X152Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444444400cc00cc)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_BLUT (
.I0(CLBLM_R_X97Y119_SLICE_X152Y119_DO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_L_X98Y120_SLICE_X154Y120_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y119_SLICE_X152Y119_BO5),
.O6(CLBLM_R_X97Y119_SLICE_X152Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y119_SLICE_X152Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y119_SLICE_X152Y119_A5Q),
.I2(CLBLL_L_X100Y122_SLICE_X156Y122_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y119_SLICE_X152Y119_AO5),
.O6(CLBLM_R_X97Y119_SLICE_X152Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X153Y119_AO5),
.Q(CLBLM_R_X97Y119_SLICE_X153Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X153Y119_CO5),
.Q(CLBLM_R_X97Y119_SLICE_X153Y119_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X153Y119_AO6),
.Q(CLBLM_R_X97Y119_SLICE_X153Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X153Y119_BO6),
.Q(CLBLM_R_X97Y119_SLICE_X153Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y119_SLICE_X153Y119_CO6),
.Q(CLBLM_R_X97Y119_SLICE_X153Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_DLUT (
.I0(CLBLM_R_X97Y119_SLICE_X153Y119_C5Q),
.I1(CLBLM_R_X97Y119_SLICE_X153Y119_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(1'b1),
.I4(CLBLM_R_X95Y119_SLICE_X150Y119_B5Q),
.I5(CLBLM_R_X97Y120_SLICE_X153Y120_BQ),
.O5(CLBLM_R_X97Y119_SLICE_X153Y119_DO5),
.O6(CLBLM_R_X97Y119_SLICE_X153Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y119_SLICE_X153Y119_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y120_SLICE_X153Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y119_SLICE_X153Y119_CO5),
.O6(CLBLM_R_X97Y119_SLICE_X153Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8aaa80aa8a008000)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y119_SLICE_X153Y119_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X97Y118_SLICE_X153Y118_AO6),
.I5(CLBLM_L_X90Y119_SLICE_X142Y119_DO6),
.O5(CLBLM_R_X97Y119_SLICE_X153Y119_BO5),
.O6(CLBLM_R_X97Y119_SLICE_X153Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X97Y119_SLICE_X153Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y119_SLICE_X153Y119_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y119_SLICE_X154Y119_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y119_SLICE_X153Y119_AO5),
.O6(CLBLM_R_X97Y119_SLICE_X153Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X152Y120_AO5),
.Q(CLBLM_R_X97Y120_SLICE_X152Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X152Y120_AO6),
.Q(CLBLM_R_X97Y120_SLICE_X152Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X152Y120_BO6),
.Q(CLBLM_R_X97Y120_SLICE_X152Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cce2e233ffe2e2)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_DLUT (
.I0(CLBLM_L_X98Y120_SLICE_X155Y120_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X97Y119_SLICE_X153Y119_DO6),
.I3(CLBLM_R_X97Y120_SLICE_X152Y120_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y119_SLICE_X150Y119_A5Q),
.O5(CLBLM_R_X97Y120_SLICE_X152Y120_DO5),
.O6(CLBLM_R_X97Y120_SLICE_X152Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3535fff035350f00)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_CLUT (
.I0(CLBLM_L_X94Y119_SLICE_X149Y119_A5Q),
.I1(CLBLM_R_X97Y120_SLICE_X152Y120_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X98Y124_SLICE_X154Y124_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X95Y119_SLICE_X150Y119_DO6),
.O5(CLBLM_R_X97Y120_SLICE_X152Y120_CO5),
.O6(CLBLM_R_X97Y120_SLICE_X152Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a00a0a0a0a)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y123_SLICE_X152Y123_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X98Y120_SLICE_X154Y120_A5Q),
.O5(CLBLM_R_X97Y120_SLICE_X152Y120_BO5),
.O6(CLBLM_R_X97Y120_SLICE_X152Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X97Y120_SLICE_X152Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y120_SLICE_X152Y120_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X97Y119_SLICE_X152Y119_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y120_SLICE_X152Y120_AO5),
.O6(CLBLM_R_X97Y120_SLICE_X152Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_AO5),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_BO5),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_CO5),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_DO5),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_AO6),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_BO6),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_CO6),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y120_SLICE_X153Y120_DO6),
.Q(CLBLM_R_X97Y120_SLICE_X153Y120_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc330000a5a50000)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_DLUT (
.I0(CLBLL_L_X102Y121_SLICE_X160Y121_AQ),
.I1(CLBLM_R_X97Y120_SLICE_X153Y120_CQ),
.I2(CLBLM_R_X97Y120_SLICE_X153Y120_DQ),
.I3(CLBLM_R_X101Y120_SLICE_X158Y120_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y120_SLICE_X153Y120_DO5),
.O6(CLBLM_R_X97Y120_SLICE_X153Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0303060906090)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_CLUT (
.I0(CLBLL_L_X100Y120_SLICE_X157Y120_BQ),
.I1(CLBLL_L_X100Y118_SLICE_X157Y118_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y121_SLICE_X153Y121_CQ),
.I4(CLBLL_L_X100Y119_SLICE_X157Y119_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y120_SLICE_X153Y120_CO5),
.O6(CLBLM_R_X97Y120_SLICE_X153Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y120_SLICE_X155Y120_A5Q),
.I2(CLBLL_L_X102Y121_SLICE_X161Y121_C5Q),
.I3(CLBLM_R_X97Y120_SLICE_X152Y120_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y120_SLICE_X153Y120_BO5),
.O6(CLBLM_R_X97Y120_SLICE_X153Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc84848484)
  ) CLBLM_R_X97Y120_SLICE_X153Y120_ALUT (
.I0(CLBLM_R_X97Y120_SLICE_X153Y120_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_L_X98Y120_SLICE_X155Y120_B5Q),
.I3(CLBLM_R_X97Y120_SLICE_X152Y120_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y120_SLICE_X153Y120_AO5),
.O6(CLBLM_R_X97Y120_SLICE_X153Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X152Y121_AO5),
.Q(CLBLM_R_X97Y121_SLICE_X152Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X152Y121_BO5),
.Q(CLBLM_R_X97Y121_SLICE_X152Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X152Y121_CO5),
.Q(CLBLM_R_X97Y121_SLICE_X152Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X152Y121_AO6),
.Q(CLBLM_R_X97Y121_SLICE_X152Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X152Y121_BO6),
.Q(CLBLM_R_X97Y121_SLICE_X152Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X152Y121_CO6),
.Q(CLBLM_R_X97Y121_SLICE_X152Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_DLUT (
.I0(CLBLM_R_X97Y121_SLICE_X152Y121_C5Q),
.I1(CLBLM_R_X97Y121_SLICE_X152Y121_CQ),
.I2(CLBLM_R_X97Y122_SLICE_X152Y122_DQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X97Y121_SLICE_X152Y121_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X152Y121_DO5),
.O6(CLBLM_R_X97Y121_SLICE_X152Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000c0c0c0c0)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y121_SLICE_X152Y121_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X97Y122_SLICE_X152Y122_DQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X152Y121_CO5),
.O6(CLBLM_R_X97Y121_SLICE_X152Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y121_SLICE_X152Y121_AQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y121_SLICE_X152Y121_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X152Y121_BO5),
.O6(CLBLM_R_X97Y121_SLICE_X152Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222aa0000aa)
  ) CLBLM_R_X97Y121_SLICE_X152Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y121_SLICE_X150Y121_BO6),
.I2(1'b1),
.I3(CLBLM_R_X97Y122_SLICE_X152Y122_D5Q),
.I4(CLBLM_R_X97Y122_SLICE_X153Y122_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X152Y121_AO5),
.O6(CLBLM_R_X97Y121_SLICE_X152Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X153Y121_AO5),
.Q(CLBLM_R_X97Y121_SLICE_X153Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X153Y121_BO5),
.Q(CLBLM_R_X97Y121_SLICE_X153Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X153Y121_CO5),
.Q(CLBLM_R_X97Y121_SLICE_X153Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X153Y121_AO6),
.Q(CLBLM_R_X97Y121_SLICE_X153Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X153Y121_BO6),
.Q(CLBLM_R_X97Y121_SLICE_X153Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y121_SLICE_X153Y121_CO6),
.Q(CLBLM_R_X97Y121_SLICE_X153Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11dd11ddf3f3c0c0)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_DLUT (
.I0(CLBLM_L_X94Y120_SLICE_X149Y120_B5Q),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X95Y121_SLICE_X151Y121_DO6),
.I3(CLBLM_R_X97Y121_SLICE_X153Y121_A5Q),
.I4(CLBLM_R_X97Y123_SLICE_X153Y123_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X97Y121_SLICE_X153Y121_DO5),
.O6(CLBLM_R_X97Y121_SLICE_X153Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_CLUT (
.I0(CLBLM_R_X97Y120_SLICE_X153Y120_C5Q),
.I1(CLBLM_L_X98Y121_SLICE_X155Y121_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X100Y121_SLICE_X157Y121_AQ),
.I4(CLBLM_R_X97Y120_SLICE_X153Y120_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X153Y121_CO5),
.O6(CLBLM_R_X97Y121_SLICE_X153Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaa00aa00a)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y124_SLICE_X154Y124_A5Q),
.I3(CLBLM_R_X97Y120_SLICE_X153Y120_A5Q),
.I4(CLBLM_R_X97Y121_SLICE_X153Y121_DO6),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X153Y121_BO5),
.O6(CLBLM_R_X97Y121_SLICE_X153Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X97Y121_SLICE_X153Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y120_SLICE_X152Y120_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X97Y121_SLICE_X153Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y121_SLICE_X153Y121_AO5),
.O6(CLBLM_R_X97Y121_SLICE_X153Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X152Y122_AO5),
.Q(CLBLM_R_X97Y122_SLICE_X152Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X152Y122_DO5),
.Q(CLBLM_R_X97Y122_SLICE_X152Y122_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X152Y122_AO6),
.Q(CLBLM_R_X97Y122_SLICE_X152Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X152Y122_BO6),
.Q(CLBLM_R_X97Y122_SLICE_X152Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X152Y122_CO6),
.Q(CLBLM_R_X97Y122_SLICE_X152Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X152Y122_DO6),
.Q(CLBLM_R_X97Y122_SLICE_X152Y122_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000f00f0000)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_DLUT (
.I0(CLBLM_R_X95Y121_SLICE_X150Y121_CO6),
.I1(1'b1),
.I2(CLBLM_R_X97Y122_SLICE_X153Y122_B5Q),
.I3(CLBLM_R_X95Y122_SLICE_X150Y122_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y122_SLICE_X152Y122_DO5),
.O6(CLBLM_R_X97Y122_SLICE_X152Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0f080c0b0308000)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_CLUT (
.I0(CLBLM_L_X98Y122_SLICE_X154Y122_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X93Y123_SLICE_X146Y123_CO6),
.I5(CLBLM_R_X97Y122_SLICE_X153Y122_AO6),
.O5(CLBLM_R_X97Y122_SLICE_X152Y122_CO5),
.O6(CLBLM_R_X97Y122_SLICE_X152Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa000a088888888)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X93Y122_SLICE_X146Y122_BO6),
.I2(CLBLM_L_X98Y121_SLICE_X154Y121_BO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y122_SLICE_X152Y122_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y122_SLICE_X152Y122_BO5),
.O6(CLBLM_R_X97Y122_SLICE_X152Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X97Y122_SLICE_X152Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y122_SLICE_X152Y122_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X98Y122_SLICE_X154Y122_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y122_SLICE_X152Y122_AO5),
.O6(CLBLM_R_X97Y122_SLICE_X152Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X153Y122_BO5),
.Q(CLBLM_R_X97Y122_SLICE_X153Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X153Y122_CO5),
.Q(CLBLM_R_X97Y122_SLICE_X153Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X153Y122_AO5),
.Q(CLBLM_R_X97Y122_SLICE_X153Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X153Y122_BO6),
.Q(CLBLM_R_X97Y122_SLICE_X153Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y122_SLICE_X153Y122_CO6),
.Q(CLBLM_R_X97Y122_SLICE_X153Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_DLUT (
.I0(CLBLM_R_X97Y122_SLICE_X153Y122_C5Q),
.I1(CLBLM_R_X97Y122_SLICE_X153Y122_CQ),
.I2(CLBLL_L_X100Y123_SLICE_X156Y123_AQ),
.I3(CLBLM_R_X97Y122_SLICE_X153Y122_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y122_SLICE_X153Y122_DO5),
.O6(CLBLM_R_X97Y122_SLICE_X153Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y122_SLICE_X153Y122_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y122_SLICE_X153Y122_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y122_SLICE_X153Y122_CO5),
.O6(CLBLM_R_X97Y122_SLICE_X153Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y122_SLICE_X155Y122_B5Q),
.I3(CLBLL_L_X100Y123_SLICE_X156Y123_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y122_SLICE_X153Y122_BO5),
.O6(CLBLM_R_X97Y122_SLICE_X153Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caa00aa00)
  ) CLBLM_R_X97Y122_SLICE_X153Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y123_SLICE_X154Y123_CQ),
.I2(CLBLM_R_X97Y122_SLICE_X153Y122_AQ),
.I3(CLBLM_L_X98Y122_SLICE_X154Y122_B5Q),
.I4(CLBLM_R_X97Y122_SLICE_X152Y122_CQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y122_SLICE_X153Y122_AO5),
.O6(CLBLM_R_X97Y122_SLICE_X153Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X152Y123_AO5),
.Q(CLBLM_R_X97Y123_SLICE_X152Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X152Y123_BO5),
.Q(CLBLM_R_X97Y123_SLICE_X152Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X152Y123_CO5),
.Q(CLBLM_R_X97Y123_SLICE_X152Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X152Y123_AO6),
.Q(CLBLM_R_X97Y123_SLICE_X152Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X152Y123_BO6),
.Q(CLBLM_R_X97Y123_SLICE_X152Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X152Y123_CO6),
.Q(CLBLM_R_X97Y123_SLICE_X152Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_DLUT (
.I0(CLBLM_L_X98Y125_SLICE_X154Y125_AQ),
.I1(CLBLM_R_X97Y124_SLICE_X152Y124_BQ),
.I2(1'b1),
.I3(CLBLM_R_X97Y123_SLICE_X152Y123_BQ),
.I4(CLBLM_R_X97Y123_SLICE_X152Y123_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y123_SLICE_X152Y123_DO5),
.O6(CLBLM_R_X97Y123_SLICE_X152Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05050c030c030)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_CLUT (
.I0(CLBLM_R_X97Y122_SLICE_X153Y122_AQ),
.I1(CLBLM_R_X97Y123_SLICE_X152Y123_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_L_X98Y121_SLICE_X154Y121_BQ),
.I4(CLBLM_R_X97Y123_SLICE_X153Y123_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y123_SLICE_X152Y123_CO5),
.O6(CLBLM_R_X97Y123_SLICE_X152Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y123_SLICE_X152Y123_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X97Y124_SLICE_X152Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y123_SLICE_X152Y123_BO5),
.O6(CLBLM_R_X97Y123_SLICE_X152Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaa00aa00a)
  ) CLBLM_R_X97Y123_SLICE_X152Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y123_SLICE_X153Y123_A5Q),
.I3(CLBLM_R_X97Y125_SLICE_X153Y125_A5Q),
.I4(CLBLM_R_X95Y123_SLICE_X151Y123_CO6),
.I5(1'b1),
.O5(CLBLM_R_X97Y123_SLICE_X152Y123_AO5),
.O6(CLBLM_R_X97Y123_SLICE_X152Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X153Y123_AO5),
.Q(CLBLM_R_X97Y123_SLICE_X153Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X153Y123_BO5),
.Q(CLBLM_R_X97Y123_SLICE_X153Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X153Y123_CO5),
.Q(CLBLM_R_X97Y123_SLICE_X153Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X153Y123_AO6),
.Q(CLBLM_R_X97Y123_SLICE_X153Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X153Y123_BO6),
.Q(CLBLM_R_X97Y123_SLICE_X153Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y123_SLICE_X153Y123_CO6),
.Q(CLBLM_R_X97Y123_SLICE_X153Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_DLUT (
.I0(CLBLM_L_X98Y124_SLICE_X154Y124_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X97Y123_SLICE_X153Y123_BQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y123_SLICE_X153Y123_B5Q),
.I5(CLBLL_L_X100Y124_SLICE_X157Y124_BQ),
.O5(CLBLM_R_X97Y123_SLICE_X153Y123_DO5),
.O6(CLBLM_R_X97Y123_SLICE_X153Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00000f090909090)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_CLUT (
.I0(CLBLM_L_X98Y123_SLICE_X154Y123_A5Q),
.I1(CLBLM_R_X97Y123_SLICE_X153Y123_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y121_SLICE_X153Y121_C5Q),
.I4(CLBLM_L_X98Y123_SLICE_X155Y123_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y123_SLICE_X153Y123_CO5),
.O6(CLBLM_R_X97Y123_SLICE_X153Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y123_SLICE_X153Y123_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X98Y124_SLICE_X154Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y123_SLICE_X153Y123_BO5),
.O6(CLBLM_R_X97Y123_SLICE_X153Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222aa0000aa)
  ) CLBLM_R_X97Y123_SLICE_X153Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y122_SLICE_X151Y122_AO6),
.I2(1'b1),
.I3(CLBLM_R_X97Y121_SLICE_X153Y121_B5Q),
.I4(CLBLM_R_X97Y123_SLICE_X153Y123_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y123_SLICE_X153Y123_AO5),
.O6(CLBLM_R_X97Y123_SLICE_X153Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y124_SLICE_X152Y124_AO5),
.Q(CLBLM_R_X97Y124_SLICE_X152Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y124_SLICE_X152Y124_BO5),
.Q(CLBLM_R_X97Y124_SLICE_X152Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y124_SLICE_X152Y124_AO6),
.Q(CLBLM_R_X97Y124_SLICE_X152Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y124_SLICE_X152Y124_BO6),
.Q(CLBLM_R_X97Y124_SLICE_X152Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y124_SLICE_X152Y124_DO5),
.O6(CLBLM_R_X97Y124_SLICE_X152Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555cccc0f0fff00)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_CLUT (
.I0(CLBLM_R_X97Y124_SLICE_X152Y124_A5Q),
.I1(CLBLM_L_X94Y124_SLICE_X149Y124_CO6),
.I2(CLBLM_R_X95Y124_SLICE_X150Y124_B5Q),
.I3(CLBLM_L_X98Y127_SLICE_X155Y127_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y124_SLICE_X152Y124_CO5),
.O6(CLBLM_R_X97Y124_SLICE_X152Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_L_X98Y125_SLICE_X154Y125_AQ),
.I3(CLBLM_R_X95Y124_SLICE_X151Y124_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y124_SLICE_X152Y124_BO5),
.O6(CLBLM_R_X97Y124_SLICE_X152Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y124_SLICE_X152Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y124_SLICE_X152Y124_A5Q),
.I2(CLBLM_R_X95Y125_SLICE_X150Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y124_SLICE_X152Y124_AO5),
.O6(CLBLM_R_X97Y124_SLICE_X152Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y124_SLICE_X153Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y124_SLICE_X153Y124_DO5),
.O6(CLBLM_R_X97Y124_SLICE_X153Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y124_SLICE_X153Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y124_SLICE_X153Y124_CO5),
.O6(CLBLM_R_X97Y124_SLICE_X153Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y124_SLICE_X153Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y124_SLICE_X153Y124_BO5),
.O6(CLBLM_R_X97Y124_SLICE_X153Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0cfa0c0afcfafc)
  ) CLBLM_R_X97Y124_SLICE_X153Y124_ALUT (
.I0(CLBLM_R_X97Y123_SLICE_X152Y123_DO6),
.I1(CLBLM_R_X101Y124_SLICE_X158Y124_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X97Y124_SLICE_X152Y124_AQ),
.I5(CLBLM_R_X95Y122_SLICE_X150Y122_A5Q),
.O5(CLBLM_R_X97Y124_SLICE_X153Y124_AO5),
.O6(CLBLM_R_X97Y124_SLICE_X153Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X152Y125_AO5),
.Q(CLBLM_R_X97Y125_SLICE_X152Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X152Y125_BO5),
.Q(CLBLM_R_X97Y125_SLICE_X152Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X152Y125_AO6),
.Q(CLBLM_R_X97Y125_SLICE_X152Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X152Y125_BO6),
.Q(CLBLM_R_X97Y125_SLICE_X152Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y125_SLICE_X152Y125_DO5),
.O6(CLBLM_R_X97Y125_SLICE_X152Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y125_SLICE_X153Y125_A5Q),
.I2(CLBLM_R_X97Y125_SLICE_X152Y125_BQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y125_SLICE_X152Y125_B5Q),
.I5(CLBLM_L_X98Y125_SLICE_X154Y125_CQ),
.O5(CLBLM_R_X97Y125_SLICE_X152Y125_CO5),
.O6(CLBLM_R_X97Y125_SLICE_X152Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y125_SLICE_X152Y125_BQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y125_SLICE_X154Y125_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y125_SLICE_X152Y125_BO5),
.O6(CLBLM_R_X97Y125_SLICE_X152Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a00aa00a)
  ) CLBLM_R_X97Y125_SLICE_X152Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y125_SLICE_X151Y125_BO6),
.I2(CLBLM_R_X97Y125_SLICE_X153Y125_B5Q),
.I3(CLBLM_R_X97Y123_SLICE_X152Y123_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y125_SLICE_X152Y125_AO5),
.O6(CLBLM_R_X97Y125_SLICE_X152Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X153Y125_AO5),
.Q(CLBLM_R_X97Y125_SLICE_X153Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X153Y125_BO5),
.Q(CLBLM_R_X97Y125_SLICE_X153Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X153Y125_AO6),
.Q(CLBLM_R_X97Y125_SLICE_X153Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y125_SLICE_X153Y125_BO6),
.Q(CLBLM_R_X97Y125_SLICE_X153Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_R_X97Y125_SLICE_X153Y125_BQ),
.I3(CLBLM_R_X97Y125_SLICE_X153Y125_AQ),
.I4(CLBLM_R_X97Y125_SLICE_X153Y125_B5Q),
.I5(CLBLM_L_X98Y126_SLICE_X154Y126_BQ),
.O5(CLBLM_R_X97Y125_SLICE_X153Y125_DO5),
.O6(CLBLM_R_X97Y125_SLICE_X153Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055d8d8aaffd8d8)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y125_SLICE_X152Y125_CO6),
.I2(CLBLL_L_X100Y126_SLICE_X156Y126_CO6),
.I3(CLBLM_R_X97Y123_SLICE_X152Y123_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_L_X98Y125_SLICE_X154Y125_B5Q),
.O5(CLBLM_R_X97Y125_SLICE_X153Y125_CO5),
.O6(CLBLM_R_X97Y125_SLICE_X153Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y125_SLICE_X153Y125_BQ),
.I2(CLBLM_R_X97Y125_SLICE_X153Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y125_SLICE_X153Y125_BO5),
.O6(CLBLM_R_X97Y125_SLICE_X153Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y125_SLICE_X153Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y126_SLICE_X154Y126_BQ),
.I2(CLBLM_R_X97Y125_SLICE_X152Y125_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y125_SLICE_X153Y125_AO5),
.O6(CLBLM_R_X97Y125_SLICE_X153Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X152Y126_AO5),
.Q(CLBLM_R_X97Y126_SLICE_X152Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X152Y126_BO5),
.Q(CLBLM_R_X97Y126_SLICE_X152Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X152Y126_AO6),
.Q(CLBLM_R_X97Y126_SLICE_X152Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X152Y126_BO6),
.Q(CLBLM_R_X97Y126_SLICE_X152Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y126_SLICE_X152Y126_DO5),
.O6(CLBLM_R_X97Y126_SLICE_X152Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X97Y127_SLICE_X152Y127_A5Q),
.I2(CLBLM_R_X97Y126_SLICE_X152Y126_BQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y126_SLICE_X152Y126_B5Q),
.I5(CLBLM_L_X98Y127_SLICE_X154Y127_BQ),
.O5(CLBLM_R_X97Y126_SLICE_X152Y126_CO5),
.O6(CLBLM_R_X97Y126_SLICE_X152Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y126_SLICE_X152Y126_BQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y127_SLICE_X154Y127_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y126_SLICE_X152Y126_BO5),
.O6(CLBLM_R_X97Y126_SLICE_X152Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa82828282)
  ) CLBLM_R_X97Y126_SLICE_X152Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y127_SLICE_X152Y127_A5Q),
.I2(CLBLM_R_X97Y125_SLICE_X152Y125_A5Q),
.I3(CLBLM_R_X95Y126_SLICE_X151Y126_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y126_SLICE_X152Y126_AO5),
.O6(CLBLM_R_X97Y126_SLICE_X152Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X153Y126_BO5),
.Q(CLBLM_R_X97Y126_SLICE_X153Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X153Y126_CO5),
.Q(CLBLM_R_X97Y126_SLICE_X153Y126_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X153Y126_AO5),
.Q(CLBLM_R_X97Y126_SLICE_X153Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X153Y126_BO6),
.Q(CLBLM_R_X97Y126_SLICE_X153Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y126_SLICE_X153Y126_CO6),
.Q(CLBLM_R_X97Y126_SLICE_X153Y126_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cacac5cac5c5ca)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_DLUT (
.I0(CLBLM_R_X97Y126_SLICE_X153Y126_BQ),
.I1(CLBLM_R_X97Y126_SLICE_X153Y126_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y126_SLICE_X153Y126_AQ),
.I4(CLBLM_R_X97Y126_SLICE_X153Y126_B5Q),
.I5(CLBLM_R_X97Y127_SLICE_X153Y127_BQ),
.O5(CLBLM_R_X97Y126_SLICE_X153Y126_DO5),
.O6(CLBLM_R_X97Y126_SLICE_X153Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50000cc330000)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_CLUT (
.I0(CLBLM_R_X97Y128_SLICE_X152Y128_AQ),
.I1(CLBLM_R_X97Y126_SLICE_X153Y126_CQ),
.I2(CLBLM_L_X94Y127_SLICE_X149Y127_B5Q),
.I3(CLBLM_L_X94Y125_SLICE_X149Y125_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y126_SLICE_X153Y126_CO5),
.O6(CLBLM_R_X97Y126_SLICE_X153Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaaa0000)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X97Y127_SLICE_X153Y127_BQ),
.I4(CLBLM_R_X97Y126_SLICE_X153Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y126_SLICE_X153Y126_BO5),
.O6(CLBLM_R_X97Y126_SLICE_X153Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_R_X97Y126_SLICE_X153Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y126_SLICE_X153Y126_BQ),
.I2(CLBLM_R_X97Y126_SLICE_X153Y126_AQ),
.I3(CLBLM_R_X97Y127_SLICE_X153Y127_BQ),
.I4(CLBLM_R_X97Y126_SLICE_X153Y126_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y126_SLICE_X153Y126_AO5),
.O6(CLBLM_R_X97Y126_SLICE_X153Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X152Y127_AO5),
.Q(CLBLM_R_X97Y127_SLICE_X152Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X152Y127_BO5),
.Q(CLBLM_R_X97Y127_SLICE_X152Y127_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X152Y127_AO6),
.Q(CLBLM_R_X97Y127_SLICE_X152Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X152Y127_BO6),
.Q(CLBLM_R_X97Y127_SLICE_X152Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_DLUT (
.I0(CLBLM_L_X98Y127_SLICE_X155Y127_AQ),
.I1(CLBLM_R_X97Y127_SLICE_X152Y127_AQ),
.I2(CLBLM_R_X97Y127_SLICE_X152Y127_BQ),
.I3(1'b1),
.I4(CLBLM_R_X97Y127_SLICE_X152Y127_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y127_SLICE_X152Y127_DO5),
.O6(CLBLM_R_X97Y127_SLICE_X152Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcc0fcc55ff5500)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_CLUT (
.I0(CLBLM_R_X95Y124_SLICE_X150Y124_C5Q),
.I1(CLBLM_R_X95Y125_SLICE_X151Y125_CO6),
.I2(CLBLM_R_X95Y126_SLICE_X151Y126_AQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_L_X98Y128_SLICE_X154Y128_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X97Y127_SLICE_X152Y127_CO5),
.O6(CLBLM_R_X97Y127_SLICE_X152Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y127_SLICE_X152Y127_BQ),
.I2(CLBLM_R_X97Y127_SLICE_X152Y127_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y127_SLICE_X152Y127_BO5),
.O6(CLBLM_R_X97Y127_SLICE_X152Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aa00aa00)
  ) CLBLM_R_X97Y127_SLICE_X152Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X97Y126_SLICE_X152Y126_B5Q),
.I4(CLBLM_L_X98Y127_SLICE_X155Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y127_SLICE_X152Y127_AO5),
.O6(CLBLM_R_X97Y127_SLICE_X152Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X153Y127_AO5),
.Q(CLBLM_R_X97Y127_SLICE_X153Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X153Y127_AO6),
.Q(CLBLM_R_X97Y127_SLICE_X153Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y127_SLICE_X153Y127_BO6),
.Q(CLBLM_R_X97Y127_SLICE_X153Y127_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y127_SLICE_X153Y127_DO5),
.O6(CLBLM_R_X97Y127_SLICE_X153Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y127_SLICE_X153Y127_CO5),
.O6(CLBLM_R_X97Y127_SLICE_X153Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heee222e200000000)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_BLUT (
.I0(CLBLM_R_X101Y127_SLICE_X159Y127_BO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X97Y126_SLICE_X153Y126_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y129_SLICE_X152Y129_AQ),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X97Y127_SLICE_X153Y127_BO5),
.O6(CLBLM_R_X97Y127_SLICE_X153Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a88228822)
  ) CLBLM_R_X97Y127_SLICE_X153Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y126_SLICE_X152Y126_A5Q),
.I2(CLBLM_R_X97Y127_SLICE_X152Y127_CO6),
.I3(CLBLM_R_X97Y127_SLICE_X152Y127_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y127_SLICE_X153Y127_AO5),
.O6(CLBLM_R_X97Y127_SLICE_X153Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y128_SLICE_X152Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y128_SLICE_X152Y128_AO6),
.Q(CLBLM_R_X97Y128_SLICE_X152Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y128_SLICE_X152Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y128_SLICE_X152Y128_DO5),
.O6(CLBLM_R_X97Y128_SLICE_X152Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y128_SLICE_X152Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y128_SLICE_X152Y128_CO5),
.O6(CLBLM_R_X97Y128_SLICE_X152Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y128_SLICE_X152Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y128_SLICE_X152Y128_BO5),
.O6(CLBLM_R_X97Y128_SLICE_X152Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2828282882828282)
  ) CLBLM_R_X97Y128_SLICE_X152Y128_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X94Y128_SLICE_X149Y128_A5Q),
.I2(CLBLM_R_X97Y129_SLICE_X152Y129_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X95Y124_SLICE_X150Y124_C5Q),
.O5(CLBLM_R_X97Y128_SLICE_X152Y128_AO5),
.O6(CLBLM_R_X97Y128_SLICE_X152Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y128_SLICE_X153Y128_BO5),
.Q(CLBLM_R_X97Y128_SLICE_X153Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y128_SLICE_X153Y128_CO5),
.Q(CLBLM_R_X97Y128_SLICE_X153Y128_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y128_SLICE_X153Y128_AO6),
.Q(CLBLM_R_X97Y128_SLICE_X153Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y128_SLICE_X153Y128_CO6),
.Q(CLBLM_R_X97Y128_SLICE_X153Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_DLUT (
.I0(CLBLM_R_X97Y128_SLICE_X153Y128_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X97Y128_SLICE_X152Y128_AQ),
.I3(CLBLM_R_X97Y128_SLICE_X153Y128_A5Q),
.I4(CLBLM_R_X97Y128_SLICE_X153Y128_AQ),
.I5(CLBLM_R_X97Y128_SLICE_X153Y128_CQ),
.O5(CLBLM_R_X97Y128_SLICE_X153Y128_DO5),
.O6(CLBLM_R_X97Y128_SLICE_X153Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y128_SLICE_X153Y128_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X97Y128_SLICE_X153Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y128_SLICE_X153Y128_CO5),
.O6(CLBLM_R_X97Y128_SLICE_X153Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y128_SLICE_X153Y128_A5Q),
.I2(CLBLM_R_X97Y128_SLICE_X153Y128_AQ),
.I3(CLBLM_R_X97Y128_SLICE_X153Y128_CQ),
.I4(CLBLM_R_X97Y128_SLICE_X153Y128_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y128_SLICE_X153Y128_BO5),
.O6(CLBLM_R_X97Y128_SLICE_X153Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacfc0c00000000)
  ) CLBLM_R_X97Y128_SLICE_X153Y128_ALUT (
.I0(CLBLM_R_X97Y129_SLICE_X152Y129_A5Q),
.I1(CLBLL_L_X102Y128_SLICE_X161Y128_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X97Y128_SLICE_X153Y128_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X97Y128_SLICE_X153Y128_AO5),
.O6(CLBLM_R_X97Y128_SLICE_X153Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y129_SLICE_X152Y129_AO5),
.Q(CLBLM_R_X97Y129_SLICE_X152Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y129_SLICE_X152Y129_BO5),
.Q(CLBLM_R_X97Y129_SLICE_X152Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y129_SLICE_X152Y129_AO6),
.Q(CLBLM_R_X97Y129_SLICE_X152Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y129_SLICE_X152Y129_BO6),
.Q(CLBLM_R_X97Y129_SLICE_X152Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y129_SLICE_X152Y129_CO6),
.Q(CLBLM_R_X97Y129_SLICE_X152Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X152Y129_DO5),
.O6(CLBLM_R_X97Y129_SLICE_X152Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a500000000)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_CLUT (
.I0(CLBLM_R_X97Y132_SLICE_X153Y132_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X95Y128_SLICE_X150Y128_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X97Y129_SLICE_X152Y129_CO5),
.O6(CLBLM_R_X97Y129_SLICE_X152Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000f0069006900)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_BLUT (
.I0(CLBLM_R_X97Y131_SLICE_X153Y131_CQ),
.I1(CLBLM_L_X94Y129_SLICE_X148Y129_AQ),
.I2(CLBLM_R_X95Y124_SLICE_X150Y124_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X95Y129_SLICE_X150Y129_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X152Y129_BO5),
.O6(CLBLM_R_X97Y129_SLICE_X152Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X97Y129_SLICE_X152Y129_ALUT (
.I0(CLBLM_L_X98Y133_SLICE_X154Y133_AQ),
.I1(CLBLM_R_X97Y129_SLICE_X152Y129_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X152Y129_AO5),
.O6(CLBLM_R_X97Y129_SLICE_X152Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y129_SLICE_X153Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X153Y129_DO5),
.O6(CLBLM_R_X97Y129_SLICE_X153Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y129_SLICE_X153Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X153Y129_CO5),
.O6(CLBLM_R_X97Y129_SLICE_X153Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y129_SLICE_X153Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X153Y129_BO5),
.O6(CLBLM_R_X97Y129_SLICE_X153Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y129_SLICE_X153Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y129_SLICE_X153Y129_AO5),
.O6(CLBLM_R_X97Y129_SLICE_X153Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y130_SLICE_X152Y130_BO5),
.Q(CLBLM_R_X97Y130_SLICE_X152Y130_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y130_SLICE_X152Y130_AO5),
.Q(CLBLM_R_X97Y130_SLICE_X152Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y130_SLICE_X152Y130_BO6),
.Q(CLBLM_R_X97Y130_SLICE_X152Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X152Y130_DO5),
.O6(CLBLM_R_X97Y130_SLICE_X152Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f099f099f066)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_CLUT (
.I0(CLBLM_R_X97Y130_SLICE_X152Y130_BQ),
.I1(CLBLM_R_X97Y130_SLICE_X152Y130_AQ),
.I2(CLBLM_R_X97Y129_SLICE_X152Y129_B5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y130_SLICE_X152Y130_B5Q),
.I5(CLBLM_L_X98Y131_SLICE_X155Y131_BQ),
.O5(CLBLM_R_X97Y130_SLICE_X152Y130_CO5),
.O6(CLBLM_R_X97Y130_SLICE_X152Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y130_SLICE_X152Y130_BQ),
.I2(1'b1),
.I3(CLBLM_L_X98Y131_SLICE_X155Y131_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X152Y130_BO5),
.O6(CLBLM_R_X97Y130_SLICE_X152Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996aaaa0000)
  ) CLBLM_R_X97Y130_SLICE_X152Y130_ALUT (
.I0(CLBLM_R_X97Y130_SLICE_X152Y130_B5Q),
.I1(CLBLM_R_X97Y130_SLICE_X152Y130_BQ),
.I2(CLBLM_R_X97Y130_SLICE_X152Y130_AQ),
.I3(CLBLM_L_X98Y131_SLICE_X155Y131_BQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X152Y130_AO5),
.O6(CLBLM_R_X97Y130_SLICE_X152Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y130_SLICE_X153Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y130_SLICE_X153Y130_AO5),
.Q(CLBLM_R_X97Y130_SLICE_X153Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y130_SLICE_X153Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y130_SLICE_X153Y130_AO6),
.Q(CLBLM_R_X97Y130_SLICE_X153Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y130_SLICE_X153Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X153Y130_DO5),
.O6(CLBLM_R_X97Y130_SLICE_X153Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y130_SLICE_X153Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X153Y130_CO5),
.O6(CLBLM_R_X97Y130_SLICE_X153Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X97Y130_SLICE_X153Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X153Y130_BO5),
.O6(CLBLM_R_X97Y130_SLICE_X153Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88228822a0a00a0a)
  ) CLBLM_R_X97Y130_SLICE_X153Y130_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y129_SLICE_X151Y129_B5Q),
.I2(CLBLM_R_X97Y130_SLICE_X153Y130_AQ),
.I3(CLBLM_R_X97Y129_SLICE_X152Y129_BQ),
.I4(CLBLM_R_X95Y130_SLICE_X151Y130_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y130_SLICE_X153Y130_AO5),
.O6(CLBLM_R_X97Y130_SLICE_X153Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X152Y131_BO5),
.Q(CLBLM_R_X97Y131_SLICE_X152Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X152Y131_AO5),
.Q(CLBLM_R_X97Y131_SLICE_X152Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X152Y131_BO6),
.Q(CLBLM_R_X97Y131_SLICE_X152Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_DLUT (
.I0(CLBLM_R_X97Y131_SLICE_X153Y131_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X97Y131_SLICE_X152Y131_AQ),
.I3(CLBLM_R_X95Y131_SLICE_X151Y131_CQ),
.I4(CLBLM_R_X97Y131_SLICE_X152Y131_B5Q),
.I5(CLBLM_R_X93Y129_SLICE_X147Y129_A5Q),
.O5(CLBLM_R_X97Y131_SLICE_X152Y131_DO5),
.O6(CLBLM_R_X97Y131_SLICE_X152Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4e4b1e4b1b1e4)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X97Y131_SLICE_X152Y131_BQ),
.I2(CLBLM_R_X93Y131_SLICE_X147Y131_AQ),
.I3(CLBLM_R_X97Y132_SLICE_X152Y132_B5Q),
.I4(CLBLM_R_X97Y132_SLICE_X152Y132_D5Q),
.I5(CLBLM_R_X97Y132_SLICE_X152Y132_BQ),
.O5(CLBLM_R_X97Y131_SLICE_X152Y131_CO5),
.O6(CLBLM_R_X97Y131_SLICE_X152Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaaa0000)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X97Y132_SLICE_X152Y132_BQ),
.I4(CLBLM_R_X95Y131_SLICE_X151Y131_CQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y131_SLICE_X152Y131_BO5),
.O6(CLBLM_R_X97Y131_SLICE_X152Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caa00aa00)
  ) CLBLM_R_X97Y131_SLICE_X152Y131_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X95Y131_SLICE_X151Y131_CQ),
.I2(CLBLM_R_X97Y131_SLICE_X152Y131_AQ),
.I3(CLBLM_R_X97Y131_SLICE_X152Y131_B5Q),
.I4(CLBLM_R_X97Y131_SLICE_X153Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y131_SLICE_X152Y131_AO5),
.O6(CLBLM_R_X97Y131_SLICE_X152Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X153Y131_BO5),
.Q(CLBLM_R_X97Y131_SLICE_X153Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X153Y131_CO5),
.Q(CLBLM_R_X97Y131_SLICE_X153Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X153Y131_AO6),
.Q(CLBLM_R_X97Y131_SLICE_X153Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X153Y131_BO6),
.Q(CLBLM_R_X97Y131_SLICE_X153Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y131_SLICE_X153Y131_CO6),
.Q(CLBLM_R_X97Y131_SLICE_X153Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cacac5cac5c5ca)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_DLUT (
.I0(CLBLM_R_X97Y131_SLICE_X153Y131_BQ),
.I1(CLBLM_R_X97Y131_SLICE_X153Y131_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y131_SLICE_X155Y131_B5Q),
.I4(CLBLM_R_X97Y131_SLICE_X153Y131_B5Q),
.I5(CLBLM_L_X98Y132_SLICE_X155Y132_BQ),
.O5(CLBLM_R_X97Y131_SLICE_X153Y131_DO5),
.O6(CLBLM_R_X97Y131_SLICE_X153Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88448844c0c00c0c)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_CLUT (
.I0(CLBLM_R_X97Y130_SLICE_X153Y130_A5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X97Y129_SLICE_X152Y129_B5Q),
.I3(CLBLM_R_X95Y131_SLICE_X151Y131_A5Q),
.I4(CLBLM_R_X97Y131_SLICE_X152Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y131_SLICE_X153Y131_CO5),
.O6(CLBLM_R_X97Y131_SLICE_X153Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaaa0000)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X98Y132_SLICE_X155Y132_BQ),
.I4(CLBLM_R_X97Y131_SLICE_X153Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y131_SLICE_X153Y131_BO5),
.O6(CLBLM_R_X97Y131_SLICE_X153Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heee222e200000000)
  ) CLBLM_R_X97Y131_SLICE_X153Y131_ALUT (
.I0(CLBLM_R_X97Y132_SLICE_X153Y132_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X97Y131_SLICE_X152Y131_AO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X95Y131_SLICE_X150Y131_AQ),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X97Y131_SLICE_X153Y131_AO5),
.O6(CLBLM_R_X97Y131_SLICE_X153Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X152Y132_AO5),
.Q(CLBLM_R_X97Y132_SLICE_X152Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X152Y132_CO5),
.Q(CLBLM_R_X97Y132_SLICE_X152Y132_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X152Y132_DO5),
.Q(CLBLM_R_X97Y132_SLICE_X152Y132_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X152Y132_AO6),
.Q(CLBLM_R_X97Y132_SLICE_X152Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X152Y132_BO6),
.Q(CLBLM_R_X97Y132_SLICE_X152Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X152Y132_DO6),
.Q(CLBLM_R_X97Y132_SLICE_X152Y132_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_DLUT (
.I0(CLBLM_R_X97Y131_SLICE_X152Y131_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X95Y132_SLICE_X151Y132_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y132_SLICE_X152Y132_DO5),
.O6(CLBLM_R_X97Y132_SLICE_X152Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999966c0c0c0c0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_CLUT (
.I0(CLBLM_R_X97Y132_SLICE_X152Y132_BQ),
.I1(CLBLM_R_X97Y132_SLICE_X152Y132_D5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X97Y131_SLICE_X152Y131_BQ),
.I4(CLBLM_R_X97Y132_SLICE_X152Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y132_SLICE_X152Y132_CO5),
.O6(CLBLM_R_X97Y132_SLICE_X152Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a808a8a8080808)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y133_SLICE_X153Y133_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X97Y132_SLICE_X152Y132_A5Q),
.I5(CLBLM_R_X97Y132_SLICE_X152Y132_CO6),
.O5(CLBLM_R_X97Y132_SLICE_X152Y132_BO5),
.O6(CLBLM_R_X97Y132_SLICE_X152Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y132_SLICE_X152Y132_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y132_SLICE_X152Y132_A5Q),
.I2(CLBLM_R_X95Y131_SLICE_X150Y131_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y132_SLICE_X152Y132_AO5),
.O6(CLBLM_R_X97Y132_SLICE_X152Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X153Y132_AO5),
.Q(CLBLM_R_X97Y132_SLICE_X153Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X153Y132_BO5),
.Q(CLBLM_R_X97Y132_SLICE_X153Y132_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X153Y132_CO5),
.Q(CLBLM_R_X97Y132_SLICE_X153Y132_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X153Y132_AO6),
.Q(CLBLM_R_X97Y132_SLICE_X153Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X153Y132_BO6),
.Q(CLBLM_R_X97Y132_SLICE_X153Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y132_SLICE_X153Y132_CO6),
.Q(CLBLM_R_X97Y132_SLICE_X153Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_DLUT (
.I0(CLBLM_L_X98Y132_SLICE_X155Y132_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X97Y131_SLICE_X153Y131_C5Q),
.I3(CLBLM_R_X97Y132_SLICE_X153Y132_A5Q),
.I4(CLBLM_R_X97Y132_SLICE_X153Y132_AQ),
.I5(CLBLM_L_X98Y133_SLICE_X155Y133_BQ),
.O5(CLBLM_R_X97Y132_SLICE_X153Y132_DO5),
.O6(CLBLM_R_X97Y132_SLICE_X153Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05050c030c030)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_CLUT (
.I0(CLBLM_R_X95Y132_SLICE_X150Y132_AQ),
.I1(CLBLM_R_X97Y132_SLICE_X153Y132_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X95Y130_SLICE_X150Y130_A5Q),
.I4(CLBLM_R_X97Y132_SLICE_X153Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y132_SLICE_X153Y132_CO5),
.O6(CLBLM_R_X97Y132_SLICE_X153Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0000aa82828282)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y132_SLICE_X153Y132_BQ),
.I2(CLBLM_R_X95Y132_SLICE_X151Y132_B5Q),
.I3(CLBLM_R_X97Y132_SLICE_X152Y132_B5Q),
.I4(CLBLM_R_X97Y131_SLICE_X153Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y132_SLICE_X153Y132_BO5),
.O6(CLBLM_R_X97Y132_SLICE_X153Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X97Y132_SLICE_X153Y132_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y133_SLICE_X155Y133_BQ),
.I2(CLBLM_R_X97Y132_SLICE_X153Y132_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X97Y132_SLICE_X153Y132_AO5),
.O6(CLBLM_R_X97Y132_SLICE_X153Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X152Y133_BO5),
.Q(CLBLM_R_X97Y133_SLICE_X152Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X152Y133_CO5),
.Q(CLBLM_R_X97Y133_SLICE_X152Y133_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X152Y133_AO6),
.Q(CLBLM_R_X97Y133_SLICE_X152Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X152Y133_CO6),
.Q(CLBLM_R_X97Y133_SLICE_X152Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f90609f9f60906)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_DLUT (
.I0(CLBLM_R_X97Y133_SLICE_X152Y133_C5Q),
.I1(CLBLM_R_X97Y133_SLICE_X152Y133_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y133_SLICE_X152Y133_A5Q),
.I4(CLBLM_R_X97Y132_SLICE_X153Y132_C5Q),
.I5(CLBLM_R_X97Y133_SLICE_X152Y133_AQ),
.O5(CLBLM_R_X97Y133_SLICE_X152Y133_DO5),
.O6(CLBLM_R_X97Y133_SLICE_X152Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff000000)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X97Y133_SLICE_X152Y133_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X97Y133_SLICE_X152Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y133_SLICE_X152Y133_CO5),
.O6(CLBLM_R_X97Y133_SLICE_X152Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69699696ff000000)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_BLUT (
.I0(CLBLM_R_X97Y133_SLICE_X152Y133_CQ),
.I1(CLBLM_R_X97Y133_SLICE_X152Y133_A5Q),
.I2(CLBLM_R_X97Y133_SLICE_X152Y133_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X97Y133_SLICE_X152Y133_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y133_SLICE_X152Y133_BO5),
.O6(CLBLM_R_X97Y133_SLICE_X152Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cccc00000000)
  ) CLBLM_R_X97Y133_SLICE_X152Y133_ALUT (
.I0(CLBLM_L_X98Y133_SLICE_X154Y133_A5Q),
.I1(CLBLM_R_X101Y135_SLICE_X158Y135_BO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X97Y133_SLICE_X152Y133_BO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X97Y133_SLICE_X152Y133_AO5),
.O6(CLBLM_R_X97Y133_SLICE_X152Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X153Y133_BO5),
.Q(CLBLM_R_X97Y133_SLICE_X153Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X153Y133_CO5),
.Q(CLBLM_R_X97Y133_SLICE_X153Y133_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X153Y133_AO6),
.Q(CLBLM_R_X97Y133_SLICE_X153Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X97Y133_SLICE_X153Y133_CO6),
.Q(CLBLM_R_X97Y133_SLICE_X153Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_DLUT (
.I0(CLBLM_R_X97Y133_SLICE_X153Y133_C5Q),
.I1(CLBLM_R_X97Y133_SLICE_X153Y133_CQ),
.I2(CLBLM_R_X97Y132_SLICE_X153Y132_BQ),
.I3(CLBLM_R_X97Y133_SLICE_X153Y133_A5Q),
.I4(CLBLM_R_X97Y133_SLICE_X153Y133_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X97Y133_SLICE_X153Y133_DO5),
.O6(CLBLM_R_X97Y133_SLICE_X153Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X97Y133_SLICE_X153Y133_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X97Y133_SLICE_X153Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X97Y133_SLICE_X153Y133_CO5),
.O6(CLBLM_R_X97Y133_SLICE_X153Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X97Y133_SLICE_X153Y133_A5Q),
.I2(CLBLM_R_X97Y133_SLICE_X153Y133_AQ),
.I3(CLBLM_R_X97Y133_SLICE_X153Y133_CQ),
.I4(CLBLM_R_X97Y133_SLICE_X153Y133_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X97Y133_SLICE_X153Y133_BO5),
.O6(CLBLM_R_X97Y133_SLICE_X153Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8fd08000000000)
  ) CLBLM_R_X97Y133_SLICE_X153Y133_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_L_X98Y133_SLICE_X155Y133_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X97Y133_SLICE_X153Y133_BO6),
.I4(CLBLM_R_X101Y136_SLICE_X159Y136_DO6),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X97Y133_SLICE_X153Y133_AO5),
.O6(CLBLM_R_X97Y133_SLICE_X153Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y110_SLICE_X158Y110_AO5),
.Q(CLBLM_R_X101Y110_SLICE_X158Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y110_SLICE_X158Y110_BO5),
.Q(CLBLM_R_X101Y110_SLICE_X158Y110_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y110_SLICE_X158Y110_AO6),
.Q(CLBLM_R_X101Y110_SLICE_X158Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y110_SLICE_X158Y110_BO6),
.Q(CLBLM_R_X101Y110_SLICE_X158Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X158Y110_DO5),
.O6(CLBLM_R_X101Y110_SLICE_X158Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_CLUT (
.I0(CLBLM_R_X101Y110_SLICE_X158Y110_BQ),
.I1(CLBLL_L_X100Y111_SLICE_X157Y111_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y110_SLICE_X158Y110_A5Q),
.I4(CLBLM_R_X101Y110_SLICE_X158Y110_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X158Y110_CO5),
.O6(CLBLM_R_X101Y110_SLICE_X158Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_BLUT (
.I0(CLBLL_L_X100Y111_SLICE_X157Y111_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y110_SLICE_X158Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X158Y110_BO5),
.O6(CLBLM_R_X101Y110_SLICE_X158Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000aa00aa00)
  ) CLBLM_R_X101Y110_SLICE_X158Y110_ALUT (
.I0(CLBLM_R_X101Y110_SLICE_X158Y110_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X100Y111_SLICE_X157Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X158Y110_AO5),
.O6(CLBLM_R_X101Y110_SLICE_X158Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y110_SLICE_X159Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X159Y110_DO5),
.O6(CLBLM_R_X101Y110_SLICE_X159Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y110_SLICE_X159Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X159Y110_CO5),
.O6(CLBLM_R_X101Y110_SLICE_X159Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y110_SLICE_X159Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X159Y110_BO5),
.O6(CLBLM_R_X101Y110_SLICE_X159Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y110_SLICE_X159Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y110_SLICE_X159Y110_AO5),
.O6(CLBLM_R_X101Y110_SLICE_X159Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X158Y111_AO5),
.Q(CLBLM_R_X101Y111_SLICE_X158Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X158Y111_BO5),
.Q(CLBLM_R_X101Y111_SLICE_X158Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X158Y111_AO6),
.Q(CLBLM_R_X101Y111_SLICE_X158Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X158Y111_BO6),
.Q(CLBLM_R_X101Y111_SLICE_X158Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_DLUT (
.I0(CLBLM_R_X101Y110_SLICE_X158Y110_AQ),
.I1(1'b1),
.I2(CLBLM_R_X101Y111_SLICE_X158Y111_BQ),
.I3(CLBLL_L_X100Y111_SLICE_X157Y111_BQ),
.I4(CLBLM_R_X101Y111_SLICE_X158Y111_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X101Y111_SLICE_X158Y111_DO5),
.O6(CLBLM_R_X101Y111_SLICE_X158Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444eeee50fa50fa)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y110_SLICE_X158Y110_CO6),
.I2(CLBLM_L_X98Y111_SLICE_X154Y111_CO6),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_A5Q),
.I4(CLBLL_L_X100Y111_SLICE_X157Y111_A5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X101Y111_SLICE_X158Y111_CO5),
.O6(CLBLM_R_X101Y111_SLICE_X158Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_BLUT (
.I0(CLBLM_R_X101Y111_SLICE_X158Y111_BQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y110_SLICE_X158Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y111_SLICE_X158Y111_BO5),
.O6(CLBLM_R_X101Y111_SLICE_X158Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X101Y111_SLICE_X158Y111_ALUT (
.I0(CLBLM_L_X98Y112_SLICE_X155Y112_AQ),
.I1(1'b1),
.I2(CLBLL_L_X100Y111_SLICE_X156Y111_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y111_SLICE_X158Y111_AO5),
.O6(CLBLM_R_X101Y111_SLICE_X158Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X159Y111_AO5),
.Q(CLBLM_R_X101Y111_SLICE_X159Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X159Y111_BO5),
.Q(CLBLM_R_X101Y111_SLICE_X159Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X159Y111_AO6),
.Q(CLBLM_R_X101Y111_SLICE_X159Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y111_SLICE_X159Y111_BO6),
.Q(CLBLM_R_X101Y111_SLICE_X159Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y111_SLICE_X159Y111_DO5),
.O6(CLBLM_R_X101Y111_SLICE_X159Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y111_SLICE_X159Y111_CO5),
.O6(CLBLM_R_X101Y111_SLICE_X159Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00aa005500)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_BLUT (
.I0(CLBLL_L_X102Y112_SLICE_X161Y112_A5Q),
.I1(1'b1),
.I2(CLBLL_L_X102Y111_SLICE_X161Y111_DO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y111_SLICE_X158Y111_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y111_SLICE_X159Y111_BO5),
.O6(CLBLM_R_X101Y111_SLICE_X159Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300a500a500)
  ) CLBLM_R_X101Y111_SLICE_X159Y111_ALUT (
.I0(CLBLM_R_X101Y111_SLICE_X159Y111_B5Q),
.I1(CLBLL_L_X102Y111_SLICE_X161Y111_CO6),
.I2(CLBLM_R_X101Y111_SLICE_X158Y111_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y111_SLICE_X159Y111_AO5),
.O6(CLBLM_R_X101Y111_SLICE_X159Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X158Y112_AO5),
.Q(CLBLM_R_X101Y112_SLICE_X158Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X158Y112_BO5),
.Q(CLBLM_R_X101Y112_SLICE_X158Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X158Y112_AO6),
.Q(CLBLM_R_X101Y112_SLICE_X158Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X158Y112_BO6),
.Q(CLBLM_R_X101Y112_SLICE_X158Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X158Y112_DO5),
.O6(CLBLM_R_X101Y112_SLICE_X158Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_CLUT (
.I0(CLBLM_R_X101Y111_SLICE_X158Y111_AQ),
.I1(CLBLM_R_X101Y112_SLICE_X158Y112_AQ),
.I2(CLBLM_L_X98Y112_SLICE_X155Y112_AQ),
.I3(CLBLM_R_X101Y112_SLICE_X158Y112_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X158Y112_CO5),
.O6(CLBLM_R_X101Y112_SLICE_X158Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00c300c300)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y112_SLICE_X158Y112_A5Q),
.I2(CLBLM_R_X101Y111_SLICE_X159Y111_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X158Y112_BO5),
.O6(CLBLM_R_X101Y112_SLICE_X158Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_R_X101Y112_SLICE_X158Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X101Y112_SLICE_X158Y112_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y111_SLICE_X158Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X158Y112_AO5),
.O6(CLBLM_R_X101Y112_SLICE_X158Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X159Y112_AO5),
.Q(CLBLM_R_X101Y112_SLICE_X159Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X159Y112_BO5),
.Q(CLBLM_R_X101Y112_SLICE_X159Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X159Y112_CO5),
.Q(CLBLM_R_X101Y112_SLICE_X159Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X159Y112_AO6),
.Q(CLBLM_R_X101Y112_SLICE_X159Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X159Y112_BO6),
.Q(CLBLM_R_X101Y112_SLICE_X159Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y112_SLICE_X159Y112_CO6),
.Q(CLBLM_R_X101Y112_SLICE_X159Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_DLUT (
.I0(CLBLM_R_X101Y112_SLICE_X159Y112_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLL_L_X100Y113_SLICE_X157Y113_AQ),
.I4(CLBLM_R_X101Y112_SLICE_X159Y112_B5Q),
.I5(CLBLM_R_X101Y112_SLICE_X159Y112_AQ),
.O5(CLBLM_R_X101Y112_SLICE_X159Y112_DO5),
.O6(CLBLM_R_X101Y112_SLICE_X159Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X100Y112_SLICE_X157Y112_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X159Y112_CO5),
.O6(CLBLM_R_X101Y112_SLICE_X159Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y112_SLICE_X159Y112_AQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y112_SLICE_X159Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X159Y112_BO5),
.O6(CLBLM_R_X101Y112_SLICE_X159Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X101Y112_SLICE_X159Y112_ALUT (
.I0(CLBLL_L_X100Y113_SLICE_X157Y113_AQ),
.I1(1'b1),
.I2(CLBLM_R_X101Y113_SLICE_X159Y113_C5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y112_SLICE_X159Y112_AO5),
.O6(CLBLM_R_X101Y112_SLICE_X159Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X158Y113_AO5),
.Q(CLBLM_R_X101Y113_SLICE_X158Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X158Y113_BO5),
.Q(CLBLM_R_X101Y113_SLICE_X158Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X158Y113_AO6),
.Q(CLBLM_R_X101Y113_SLICE_X158Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X158Y113_BO6),
.Q(CLBLM_R_X101Y113_SLICE_X158Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_DLUT (
.I0(CLBLM_R_X101Y113_SLICE_X158Y113_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLL_L_X100Y113_SLICE_X156Y113_CQ),
.I3(CLBLM_R_X101Y113_SLICE_X158Y113_A5Q),
.I4(CLBLM_R_X101Y113_SLICE_X158Y113_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y113_SLICE_X158Y113_DO5),
.O6(CLBLM_R_X101Y113_SLICE_X158Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h53ff530f53f05300)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_CLUT (
.I0(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I1(CLBLL_L_X102Y113_SLICE_X160Y113_A5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y113_SLICE_X158Y113_DO6),
.I5(CLBLL_L_X100Y113_SLICE_X156Y113_DO6),
.O5(CLBLM_R_X101Y113_SLICE_X158Y113_CO5),
.O6(CLBLM_R_X101Y113_SLICE_X158Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_BLUT (
.I0(CLBLL_L_X100Y113_SLICE_X156Y113_CQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y113_SLICE_X158Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y113_SLICE_X158Y113_BO5),
.O6(CLBLM_R_X101Y113_SLICE_X158Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X101Y113_SLICE_X158Y113_ALUT (
.I0(CLBLM_R_X101Y113_SLICE_X158Y113_B5Q),
.I1(CLBLL_L_X100Y114_SLICE_X156Y114_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y113_SLICE_X158Y113_AO5),
.O6(CLBLM_R_X101Y113_SLICE_X158Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X159Y113_CO5),
.Q(CLBLM_R_X101Y113_SLICE_X159Y113_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X159Y113_BO5),
.Q(CLBLM_R_X101Y113_SLICE_X159Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X159Y113_AO5),
.Q(CLBLM_R_X101Y113_SLICE_X159Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y113_SLICE_X159Y113_CO6),
.Q(CLBLM_R_X101Y113_SLICE_X159Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_DLUT (
.I0(CLBLL_L_X100Y115_SLICE_X156Y115_BQ),
.I1(CLBLM_R_X101Y113_SLICE_X159Y113_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X101Y113_SLICE_X159Y113_C5Q),
.I5(CLBLM_R_X101Y112_SLICE_X159Y112_A5Q),
.O5(CLBLM_R_X101Y113_SLICE_X159Y113_DO5),
.O6(CLBLM_R_X101Y113_SLICE_X159Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_CLUT (
.I0(CLBLL_L_X100Y115_SLICE_X156Y115_BQ),
.I1(CLBLM_R_X101Y113_SLICE_X159Y113_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y113_SLICE_X159Y113_CO5),
.O6(CLBLM_R_X101Y113_SLICE_X159Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa555555cccc0000)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_BLUT (
.I0(CLBLM_R_X101Y114_SLICE_X158Y114_DO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y113_SLICE_X159Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y113_SLICE_X159Y113_BO5),
.O6(CLBLM_R_X101Y113_SLICE_X159Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05fc0c0c0c0)
  ) CLBLM_R_X101Y113_SLICE_X159Y113_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I3(CLBLM_R_X101Y113_SLICE_X158Y113_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y113_SLICE_X159Y113_AO5),
.O6(CLBLM_R_X101Y113_SLICE_X159Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y114_SLICE_X158Y114_AO5),
.Q(CLBLM_R_X101Y114_SLICE_X158Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y114_SLICE_X158Y114_BO5),
.Q(CLBLM_R_X101Y114_SLICE_X158Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y114_SLICE_X158Y114_AO6),
.Q(CLBLM_R_X101Y114_SLICE_X158Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y114_SLICE_X158Y114_BO6),
.Q(CLBLM_R_X101Y114_SLICE_X158Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_DLUT (
.I0(CLBLM_R_X101Y113_SLICE_X158Y113_AQ),
.I1(1'b1),
.I2(CLBLM_R_X101Y114_SLICE_X158Y114_AQ),
.I3(CLBLM_R_X101Y114_SLICE_X158Y114_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X100Y114_SLICE_X156Y114_BQ),
.O5(CLBLM_R_X101Y114_SLICE_X158Y114_DO5),
.O6(CLBLM_R_X101Y114_SLICE_X158Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11fc1130ddfcdd30)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_CLUT (
.I0(CLBLM_R_X101Y114_SLICE_X158Y114_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_L_X98Y115_SLICE_X155Y115_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y114_SLICE_X158Y114_DO6),
.I5(CLBLM_R_X101Y113_SLICE_X159Y113_BQ),
.O5(CLBLM_R_X101Y114_SLICE_X158Y114_CO5),
.O6(CLBLM_R_X101Y114_SLICE_X158Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000f0099009900)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_BLUT (
.I0(CLBLM_R_X101Y118_SLICE_X159Y118_A5Q),
.I1(CLBLM_R_X101Y114_SLICE_X158Y114_BQ),
.I2(CLBLL_L_X102Y113_SLICE_X160Y113_A5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y114_SLICE_X158Y114_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y114_SLICE_X158Y114_BO5),
.O6(CLBLM_R_X101Y114_SLICE_X158Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_R_X101Y114_SLICE_X158Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X101Y114_SLICE_X158Y114_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y113_SLICE_X158Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y114_SLICE_X158Y114_AO5),
.O6(CLBLM_R_X101Y114_SLICE_X158Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y114_SLICE_X159Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y114_SLICE_X159Y114_DO5),
.O6(CLBLM_R_X101Y114_SLICE_X159Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y114_SLICE_X159Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y114_SLICE_X159Y114_CO5),
.O6(CLBLM_R_X101Y114_SLICE_X159Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y114_SLICE_X159Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y114_SLICE_X159Y114_BO5),
.O6(CLBLM_R_X101Y114_SLICE_X159Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y114_SLICE_X159Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y114_SLICE_X159Y114_AO5),
.O6(CLBLM_R_X101Y114_SLICE_X159Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y115_SLICE_X158Y115_AO5),
.Q(CLBLM_R_X101Y115_SLICE_X158Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y115_SLICE_X158Y115_BO5),
.Q(CLBLM_R_X101Y115_SLICE_X158Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y115_SLICE_X158Y115_AO6),
.Q(CLBLM_R_X101Y115_SLICE_X158Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y115_SLICE_X158Y115_BO6),
.Q(CLBLM_R_X101Y115_SLICE_X158Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X158Y115_DO5),
.O6(CLBLM_R_X101Y115_SLICE_X158Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_CLUT (
.I0(CLBLL_L_X100Y117_SLICE_X157Y117_BQ),
.I1(CLBLM_R_X101Y115_SLICE_X158Y115_AQ),
.I2(CLBLM_R_X101Y115_SLICE_X158Y115_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X101Y115_SLICE_X158Y115_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X158Y115_CO5),
.O6(CLBLM_R_X101Y115_SLICE_X158Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y115_SLICE_X158Y115_AQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y115_SLICE_X158Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X158Y115_BO5),
.O6(CLBLM_R_X101Y115_SLICE_X158Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cccc0000)
  ) CLBLM_R_X101Y115_SLICE_X158Y115_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLL_L_X100Y117_SLICE_X157Y117_BQ),
.I3(1'b1),
.I4(CLBLL_L_X100Y115_SLICE_X157Y115_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X158Y115_AO5),
.O6(CLBLM_R_X101Y115_SLICE_X158Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y115_SLICE_X159Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X159Y115_DO5),
.O6(CLBLM_R_X101Y115_SLICE_X159Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y115_SLICE_X159Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X159Y115_CO5),
.O6(CLBLM_R_X101Y115_SLICE_X159Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y115_SLICE_X159Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X159Y115_BO5),
.O6(CLBLM_R_X101Y115_SLICE_X159Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y115_SLICE_X159Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y115_SLICE_X159Y115_AO5),
.O6(CLBLM_R_X101Y115_SLICE_X159Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X158Y116_AO5),
.Q(CLBLM_R_X101Y116_SLICE_X158Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X158Y116_BO5),
.Q(CLBLM_R_X101Y116_SLICE_X158Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X158Y116_AO6),
.Q(CLBLM_R_X101Y116_SLICE_X158Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X158Y116_BO6),
.Q(CLBLM_R_X101Y116_SLICE_X158Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y116_SLICE_X158Y116_AQ),
.I2(CLBLM_R_X101Y116_SLICE_X158Y116_BQ),
.I3(CLBLL_L_X100Y115_SLICE_X156Y115_CQ),
.I4(CLBLM_R_X101Y116_SLICE_X158Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_DO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f033ff55f03300)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_CLUT (
.I0(CLBLM_R_X101Y113_SLICE_X159Y113_AQ),
.I1(CLBLM_R_X101Y114_SLICE_X158Y114_B5Q),
.I2(CLBLM_R_X101Y116_SLICE_X159Y116_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X100Y116_SLICE_X157Y116_DO6),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_CO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y116_SLICE_X158Y116_BQ),
.I2(CLBLM_R_X101Y116_SLICE_X158Y116_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_BO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y115_SLICE_X156Y115_CQ),
.I2(CLBLL_L_X100Y116_SLICE_X156Y116_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_AO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X159Y116_CO5),
.Q(CLBLM_R_X101Y116_SLICE_X159Y116_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X159Y116_CO6),
.Q(CLBLM_R_X101Y116_SLICE_X159Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_DLUT (
.I0(CLBLM_R_X101Y116_SLICE_X159Y116_C5Q),
.I1(CLBLL_L_X100Y116_SLICE_X157Y116_BQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y118_SLICE_X159Y118_A5Q),
.I4(CLBLM_R_X101Y116_SLICE_X159Y116_CQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_DO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y116_SLICE_X159Y116_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X100Y116_SLICE_X157Y116_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_CO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f00ffa0a0a0a0)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y113_SLICE_X159Y113_AQ),
.I3(CLBLM_R_X101Y116_SLICE_X159Y116_DO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_BO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3300ff88888888)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y117_SLICE_X159Y117_AQ),
.I2(1'b1),
.I3(CLBLM_R_X101Y115_SLICE_X158Y115_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_AO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X158Y117_BO5),
.Q(CLBLM_R_X101Y117_SLICE_X158Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X158Y117_AO6),
.Q(CLBLM_R_X101Y117_SLICE_X158Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X158Y117_BO6),
.Q(CLBLM_R_X101Y117_SLICE_X158Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aaffaa33f033f0)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_DLUT (
.I0(CLBLM_R_X101Y118_SLICE_X158Y118_DO6),
.I1(CLBLM_R_X101Y117_SLICE_X158Y117_AQ),
.I2(CLBLM_R_X97Y117_SLICE_X152Y117_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y117_SLICE_X161Y117_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_DO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h550fffcc550f00cc)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_CLUT (
.I0(CLBLM_R_X101Y117_SLICE_X159Y117_AQ),
.I1(CLBLL_L_X100Y118_SLICE_X156Y118_CO6),
.I2(CLBLM_R_X101Y117_SLICE_X158Y117_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X101Y115_SLICE_X158Y115_CO6),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_CO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50000cc330000)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_BLUT (
.I0(CLBLM_R_X101Y115_SLICE_X158Y115_B5Q),
.I1(CLBLM_R_X101Y117_SLICE_X158Y117_BQ),
.I2(CLBLM_R_X101Y117_SLICE_X158Y117_AQ),
.I3(CLBLL_L_X102Y116_SLICE_X161Y116_A5Q),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_BO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666999900000000)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_ALUT (
.I0(CLBLL_L_X100Y118_SLICE_X157Y118_C5Q),
.I1(CLBLM_R_X101Y117_SLICE_X159Y117_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y117_SLICE_X159Y117_CQ),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_AO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X159Y117_BO5),
.Q(CLBLM_R_X101Y117_SLICE_X159Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X159Y117_AO6),
.Q(CLBLM_R_X101Y117_SLICE_X159Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X159Y117_BO6),
.Q(CLBLM_R_X101Y117_SLICE_X159Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y117_SLICE_X159Y117_CO6),
.Q(CLBLM_R_X101Y117_SLICE_X159Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_DO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00cc00cc00cc00c)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y114_SLICE_X158Y114_B5Q),
.I3(CLBLM_R_X101Y118_SLICE_X159Y118_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_CO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y117_SLICE_X160Y117_AQ),
.I2(CLBLM_R_X101Y118_SLICE_X158Y118_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_BO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00c30fc30f)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y118_SLICE_X158Y118_DO6),
.I3(CLBLL_L_X102Y117_SLICE_X161Y117_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_AO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X158Y118_AO5),
.Q(CLBLM_R_X101Y118_SLICE_X158Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X158Y118_BO5),
.Q(CLBLM_R_X101Y118_SLICE_X158Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X158Y118_AO6),
.Q(CLBLM_R_X101Y118_SLICE_X158Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X158Y118_BO6),
.Q(CLBLM_R_X101Y118_SLICE_X158Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X158Y118_CO6),
.Q(CLBLM_R_X101Y118_SLICE_X158Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y118_SLICE_X158Y118_AQ),
.I2(CLBLM_R_X101Y117_SLICE_X159Y117_B5Q),
.I3(CLBLM_R_X101Y118_SLICE_X158Y118_BQ),
.I4(CLBLM_R_X101Y118_SLICE_X158Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_DO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6090609060906090)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_CLUT (
.I0(CLBLL_L_X102Y117_SLICE_X160Y117_B5Q),
.I1(CLBLM_R_X101Y119_SLICE_X158Y119_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y117_SLICE_X159Y117_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_CO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y118_SLICE_X158Y118_BQ),
.I2(CLBLM_R_X101Y118_SLICE_X158Y118_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_BO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa0000aaaa)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X101Y117_SLICE_X158Y117_DO6),
.I4(CLBLL_L_X100Y120_SLICE_X157Y120_DO6),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_AO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X159Y118_AO5),
.Q(CLBLM_R_X101Y118_SLICE_X159Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X159Y118_BO5),
.Q(CLBLM_R_X101Y118_SLICE_X159Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X159Y118_AO6),
.Q(CLBLM_R_X101Y118_SLICE_X159Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y118_SLICE_X159Y118_BO6),
.Q(CLBLM_R_X101Y118_SLICE_X159Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y116_SLICE_X159Y116_BO5),
.Q(CLBLM_R_X101Y118_SLICE_X159Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y118_SLICE_X159Y118_AQ),
.I2(1'b1),
.I3(CLBLM_R_X101Y118_SLICE_X159Y118_BQ),
.I4(CLBLM_R_X101Y118_SLICE_X159Y118_B5Q),
.I5(CLBLL_L_X100Y118_SLICE_X157Y118_AQ),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_DO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22fa225077fa7750)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y118_SLICE_X159Y118_CQ),
.I2(CLBLM_L_X98Y117_SLICE_X155Y117_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y118_SLICE_X159Y118_DO6),
.I5(CLBLM_R_X101Y117_SLICE_X159Y117_CQ),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_CO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y118_SLICE_X159Y118_BQ),
.I2(CLBLM_R_X101Y118_SLICE_X159Y118_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_BO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y118_SLICE_X157Y118_AQ),
.I2(CLBLM_R_X101Y116_SLICE_X159Y116_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_AO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X158Y119_AO5),
.Q(CLBLM_R_X101Y119_SLICE_X158Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X158Y119_AO6),
.Q(CLBLM_R_X101Y119_SLICE_X158Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X158Y119_BO6),
.Q(CLBLM_R_X101Y119_SLICE_X158Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X158Y119_CO6),
.Q(CLBLM_R_X101Y119_SLICE_X158Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_DO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9090909090909090)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_CLUT (
.I0(CLBLM_R_X101Y123_SLICE_X159Y123_C5Q),
.I1(CLBLM_R_X101Y119_SLICE_X159Y119_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_CO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha088aaaaa0880000)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y119_SLICE_X159Y119_DO6),
.I2(CLBLL_L_X102Y117_SLICE_X161Y117_CQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X98Y119_SLICE_X154Y119_DO6),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_BO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLL_L_X100Y119_SLICE_X157Y119_CQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y120_SLICE_X158Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_AO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X159Y119_AO5),
.Q(CLBLM_R_X101Y119_SLICE_X159Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X159Y119_BO5),
.Q(CLBLM_R_X101Y119_SLICE_X159Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X159Y119_AO6),
.Q(CLBLM_R_X101Y119_SLICE_X159Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y119_SLICE_X159Y119_BO6),
.Q(CLBLM_R_X101Y119_SLICE_X159Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y119_SLICE_X159Y119_BQ),
.I3(CLBLM_R_X101Y119_SLICE_X159Y119_AQ),
.I4(CLBLM_R_X101Y119_SLICE_X159Y119_B5Q),
.I5(CLBLM_R_X101Y119_SLICE_X158Y119_BQ),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_DO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_CLUT (
.I0(CLBLL_L_X102Y117_SLICE_X161Y117_CQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y119_SLICE_X159Y119_BQ),
.I3(CLBLM_R_X101Y119_SLICE_X159Y119_AQ),
.I4(CLBLM_R_X101Y119_SLICE_X159Y119_B5Q),
.I5(CLBLM_R_X101Y119_SLICE_X158Y119_BQ),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_CO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y119_SLICE_X159Y119_BQ),
.I2(CLBLM_R_X101Y119_SLICE_X159Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_BO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y120_SLICE_X159Y120_B5Q),
.I3(CLBLM_R_X101Y119_SLICE_X158Y119_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_AO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X158Y120_BO5),
.Q(CLBLM_R_X101Y120_SLICE_X158Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X158Y120_CO5),
.Q(CLBLM_R_X101Y120_SLICE_X158Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X158Y120_AO6),
.Q(CLBLM_R_X101Y120_SLICE_X158Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X158Y120_CO6),
.Q(CLBLM_R_X101Y120_SLICE_X158Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeededde12212112)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_DLUT (
.I0(CLBLM_R_X101Y120_SLICE_X158Y120_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y120_SLICE_X158Y120_AQ),
.I3(CLBLM_R_X101Y120_SLICE_X158Y120_A5Q),
.I4(CLBLM_R_X101Y119_SLICE_X158Y119_AQ),
.I5(CLBLL_L_X102Y120_SLICE_X160Y120_CQ),
.O5(CLBLM_R_X101Y120_SLICE_X158Y120_DO5),
.O6(CLBLM_R_X101Y120_SLICE_X158Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000a0a0a0a0)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_CLUT (
.I0(CLBLM_R_X101Y119_SLICE_X158Y119_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLL_L_X100Y121_SLICE_X157Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y120_SLICE_X158Y120_CO5),
.O6(CLBLM_R_X101Y120_SLICE_X158Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33caaaa0000)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y120_SLICE_X158Y120_A5Q),
.I2(CLBLM_R_X101Y119_SLICE_X158Y119_AQ),
.I3(CLBLM_R_X101Y120_SLICE_X158Y120_AQ),
.I4(CLBLM_R_X101Y120_SLICE_X158Y120_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y120_SLICE_X158Y120_BO5),
.O6(CLBLM_R_X101Y120_SLICE_X158Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a28080aa228800)
  ) CLBLM_R_X101Y120_SLICE_X158Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLL_L_X100Y120_SLICE_X157Y120_A5Q),
.I3(CLBLM_R_X101Y120_SLICE_X158Y120_BO6),
.I4(CLBLM_L_X94Y121_SLICE_X148Y121_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y120_SLICE_X158Y120_AO5),
.O6(CLBLM_R_X101Y120_SLICE_X158Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X159Y120_BO5),
.Q(CLBLM_R_X101Y120_SLICE_X159Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X159Y120_AO6),
.Q(CLBLM_R_X101Y120_SLICE_X159Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y120_SLICE_X159Y120_BO6),
.Q(CLBLM_R_X101Y120_SLICE_X159Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966669966999966)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_DLUT (
.I0(CLBLM_R_X101Y120_SLICE_X159Y120_BQ),
.I1(CLBLM_R_X101Y120_SLICE_X159Y120_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y120_SLICE_X159Y120_B5Q),
.I5(CLBLM_R_X101Y119_SLICE_X159Y119_A5Q),
.O5(CLBLM_R_X101Y120_SLICE_X159Y120_DO5),
.O6(CLBLM_R_X101Y120_SLICE_X159Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696696996)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_CLUT (
.I0(CLBLM_R_X101Y119_SLICE_X159Y119_A5Q),
.I1(CLBLM_R_X101Y120_SLICE_X159Y120_AQ),
.I2(CLBLM_R_X101Y120_SLICE_X159Y120_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y120_SLICE_X159Y120_B5Q),
.I5(CLBLL_L_X102Y122_SLICE_X160Y122_BQ),
.O5(CLBLM_R_X101Y120_SLICE_X159Y120_CO5),
.O6(CLBLM_R_X101Y120_SLICE_X159Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y120_SLICE_X159Y120_BQ),
.I2(CLBLM_R_X101Y120_SLICE_X159Y120_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y120_SLICE_X159Y120_BO5),
.O6(CLBLM_R_X101Y120_SLICE_X159Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacaff0000000000)
  ) CLBLM_R_X101Y120_SLICE_X159Y120_ALUT (
.I0(CLBLM_R_X101Y120_SLICE_X159Y120_DO6),
.I1(CLBLL_L_X102Y122_SLICE_X160Y122_BQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_L_X98Y120_SLICE_X155Y120_CO6),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y120_SLICE_X159Y120_AO5),
.O6(CLBLM_R_X101Y120_SLICE_X159Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X158Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X158Y121_AO5),
.Q(CLBLM_R_X101Y121_SLICE_X158Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X158Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X158Y121_AO6),
.Q(CLBLM_R_X101Y121_SLICE_X158Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y121_SLICE_X158Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y121_SLICE_X158Y121_DO5),
.O6(CLBLM_R_X101Y121_SLICE_X158Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X101Y121_SLICE_X158Y121_CLUT (
.I0(CLBLL_L_X100Y122_SLICE_X157Y122_AQ),
.I1(CLBLM_R_X101Y121_SLICE_X158Y121_AQ),
.I2(CLBLM_R_X101Y121_SLICE_X159Y121_B5Q),
.I3(CLBLM_R_X101Y121_SLICE_X158Y121_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X101Y121_SLICE_X158Y121_CO5),
.O6(CLBLM_R_X101Y121_SLICE_X158Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500ffccccf0f0)
  ) CLBLM_R_X101Y121_SLICE_X158Y121_BLUT (
.I0(CLBLL_L_X100Y122_SLICE_X156Y122_AQ),
.I1(CLBLM_R_X101Y121_SLICE_X159Y121_DO6),
.I2(CLBLM_R_X103Y121_SLICE_X163Y121_DO6),
.I3(CLBLL_L_X100Y121_SLICE_X156Y121_C5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y121_SLICE_X158Y121_BO5),
.O6(CLBLM_R_X101Y121_SLICE_X158Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X101Y121_SLICE_X158Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y121_SLICE_X158Y121_AQ),
.I3(1'b1),
.I4(CLBLL_L_X100Y122_SLICE_X157Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y121_SLICE_X158Y121_AO5),
.O6(CLBLM_R_X101Y121_SLICE_X158Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X159Y121_AO5),
.Q(CLBLM_R_X101Y121_SLICE_X159Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X159Y121_BO5),
.Q(CLBLM_R_X101Y121_SLICE_X159Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X159Y121_CO5),
.Q(CLBLM_R_X101Y121_SLICE_X159Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X159Y121_AO6),
.Q(CLBLM_R_X101Y121_SLICE_X159Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X159Y121_BO6),
.Q(CLBLM_R_X101Y121_SLICE_X159Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y121_SLICE_X159Y121_CO6),
.Q(CLBLM_R_X101Y121_SLICE_X159Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_DLUT (
.I0(CLBLM_R_X101Y121_SLICE_X159Y121_C5Q),
.I1(CLBLM_R_X101Y121_SLICE_X159Y121_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y121_SLICE_X159Y121_BQ),
.I4(1'b1),
.I5(CLBLM_R_X101Y121_SLICE_X159Y121_AQ),
.O5(CLBLM_R_X101Y121_SLICE_X159Y121_DO5),
.O6(CLBLM_R_X101Y121_SLICE_X159Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y121_SLICE_X159Y121_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y121_SLICE_X159Y121_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y121_SLICE_X159Y121_CO5),
.O6(CLBLM_R_X101Y121_SLICE_X159Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y121_SLICE_X159Y121_AQ),
.I3(CLBLM_R_X101Y121_SLICE_X158Y121_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y121_SLICE_X159Y121_BO5),
.O6(CLBLM_R_X101Y121_SLICE_X159Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222a0a00a0a)
  ) CLBLM_R_X101Y121_SLICE_X159Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y121_SLICE_X158Y121_BO6),
.I2(CLBLM_R_X101Y122_SLICE_X159Y122_B5Q),
.I3(1'b1),
.I4(CLBLL_L_X100Y122_SLICE_X157Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y121_SLICE_X159Y121_AO5),
.O6(CLBLM_R_X101Y121_SLICE_X159Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X158Y122_AO5),
.Q(CLBLM_R_X101Y122_SLICE_X158Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X158Y122_BO5),
.Q(CLBLM_R_X101Y122_SLICE_X158Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X158Y122_AO6),
.Q(CLBLM_R_X101Y122_SLICE_X158Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X158Y122_BO6),
.Q(CLBLM_R_X101Y122_SLICE_X158Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y122_SLICE_X159Y122_A5Q),
.I2(CLBLM_R_X101Y122_SLICE_X158Y122_BQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y122_SLICE_X158Y122_B5Q),
.I5(CLBLL_L_X102Y122_SLICE_X160Y122_CQ),
.O5(CLBLM_R_X101Y122_SLICE_X158Y122_DO5),
.O6(CLBLM_R_X101Y122_SLICE_X158Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32ba76fe109854dc)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y122_SLICE_X161Y122_DO6),
.I3(CLBLM_R_X101Y122_SLICE_X158Y122_A5Q),
.I4(CLBLL_L_X100Y122_SLICE_X157Y122_A5Q),
.I5(CLBLM_R_X101Y122_SLICE_X158Y122_DO6),
.O5(CLBLM_R_X101Y122_SLICE_X158Y122_CO5),
.O6(CLBLM_R_X101Y122_SLICE_X158Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y122_SLICE_X158Y122_BQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y122_SLICE_X160Y122_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y122_SLICE_X158Y122_BO5),
.O6(CLBLM_R_X101Y122_SLICE_X158Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X101Y122_SLICE_X158Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y122_SLICE_X158Y122_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X101Y124_SLICE_X158Y124_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y122_SLICE_X158Y122_AO5),
.O6(CLBLM_R_X101Y122_SLICE_X158Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X159Y122_AO5),
.Q(CLBLM_R_X101Y122_SLICE_X159Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X159Y122_BO5),
.Q(CLBLM_R_X101Y122_SLICE_X159Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X159Y122_AO6),
.Q(CLBLM_R_X101Y122_SLICE_X159Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y122_SLICE_X159Y122_BO6),
.Q(CLBLM_R_X101Y122_SLICE_X159Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y122_SLICE_X159Y122_AQ),
.I2(CLBLM_R_X101Y122_SLICE_X159Y122_BQ),
.I3(CLBLL_L_X102Y122_SLICE_X161Y122_CQ),
.I4(CLBLM_R_X101Y122_SLICE_X159Y122_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y122_SLICE_X159Y122_DO5),
.O6(CLBLM_R_X101Y122_SLICE_X159Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff550033f033f0)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_CLUT (
.I0(CLBLM_R_X101Y122_SLICE_X158Y122_AQ),
.I1(CLBLM_R_X101Y121_SLICE_X159Y121_A5Q),
.I2(CLBLM_R_X103Y122_SLICE_X162Y122_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y122_SLICE_X159Y122_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X101Y122_SLICE_X159Y122_CO5),
.O6(CLBLM_R_X101Y122_SLICE_X159Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y122_SLICE_X159Y122_BQ),
.I2(CLBLM_R_X101Y122_SLICE_X159Y122_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y122_SLICE_X159Y122_BO5),
.O6(CLBLM_R_X101Y122_SLICE_X159Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X101Y122_SLICE_X159Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y122_SLICE_X161Y122_CQ),
.I2(1'b1),
.I3(CLBLM_R_X101Y122_SLICE_X158Y122_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y122_SLICE_X159Y122_AO5),
.O6(CLBLM_R_X101Y122_SLICE_X159Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.Q(CLBLM_R_X101Y123_SLICE_X158Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X158Y123_BO5),
.Q(CLBLM_R_X101Y123_SLICE_X158Y123_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X158Y123_AO6),
.Q(CLBLM_R_X101Y123_SLICE_X158Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X158Y123_BO6),
.Q(CLBLM_R_X101Y123_SLICE_X158Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_AQ),
.I2(CLBLM_R_X101Y123_SLICE_X158Y123_BQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y123_SLICE_X158Y123_B5Q),
.I5(CLBLL_L_X102Y123_SLICE_X161Y123_AQ),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_DO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32ba76fe109854dc)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X102Y122_SLICE_X160Y122_DO6),
.I3(CLBLM_R_X101Y124_SLICE_X158Y124_AQ),
.I4(CLBLL_L_X100Y123_SLICE_X156Y123_A5Q),
.I5(CLBLM_R_X101Y123_SLICE_X158Y123_DO6),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_CO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_BQ),
.I2(CLBLM_R_X101Y123_SLICE_X158Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_BO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y124_SLICE_X158Y124_B5Q),
.I3(CLBLL_L_X102Y123_SLICE_X161Y123_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X159Y123_AO5),
.Q(CLBLM_R_X101Y123_SLICE_X159Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X159Y123_CO5),
.Q(CLBLM_R_X101Y123_SLICE_X159Y123_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X159Y123_AO6),
.Q(CLBLM_R_X101Y123_SLICE_X159Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X159Y123_BO6),
.Q(CLBLM_R_X101Y123_SLICE_X159Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y123_SLICE_X159Y123_CO6),
.Q(CLBLM_R_X101Y123_SLICE_X159Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_DO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h90909090f00000f0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_CLUT (
.I0(CLBLL_L_X102Y124_SLICE_X160Y124_C5Q),
.I1(CLBLL_L_X102Y124_SLICE_X160Y124_D5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLL_L_X102Y123_SLICE_X160Y123_B5Q),
.I4(CLBLM_R_X101Y123_SLICE_X159Y123_CQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_CO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff5f00000f5f)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_BLUT (
.I0(CLBLL_L_X102Y122_SLICE_X160Y122_DO6),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y123_SLICE_X161Y123_BO6),
.I5(CLBLM_R_X101Y123_SLICE_X159Y123_A5Q),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_BO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000088888888)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_ALUT (
.I0(CLBLL_L_X102Y126_SLICE_X160Y126_AQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y123_SLICE_X159Y123_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_AO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y124_SLICE_X158Y124_AO5),
.Q(CLBLM_R_X101Y124_SLICE_X158Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y124_SLICE_X158Y124_BO5),
.Q(CLBLM_R_X101Y124_SLICE_X158Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y124_SLICE_X158Y124_AO6),
.Q(CLBLM_R_X101Y124_SLICE_X158Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y124_SLICE_X158Y124_BO6),
.Q(CLBLM_R_X101Y124_SLICE_X158Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y123_SLICE_X158Y123_A5Q),
.I2(CLBLM_R_X101Y124_SLICE_X159Y124_AQ),
.I3(CLBLM_R_X101Y124_SLICE_X158Y124_BQ),
.I4(CLBLM_R_X101Y124_SLICE_X158Y124_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_DO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h37bf159d26ae048c)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLL_L_X100Y123_SLICE_X156Y123_B5Q),
.I3(CLBLM_R_X101Y124_SLICE_X158Y124_A5Q),
.I4(CLBLM_R_X101Y124_SLICE_X158Y124_DO6),
.I5(CLBLL_L_X102Y125_SLICE_X161Y125_DO6),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_CO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y124_SLICE_X158Y124_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y124_SLICE_X159Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_BO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X101Y124_SLICE_X158Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y124_SLICE_X158Y124_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X100Y125_SLICE_X157Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X158Y124_AO5),
.O6(CLBLM_R_X101Y124_SLICE_X158Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y124_SLICE_X159Y124_AO5),
.Q(CLBLM_R_X101Y124_SLICE_X159Y124_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y124_SLICE_X159Y124_AO6),
.Q(CLBLM_R_X101Y124_SLICE_X159Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_DO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_CO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_BO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a22888822)
  ) CLBLM_R_X101Y124_SLICE_X159Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_C5Q),
.I2(CLBLM_R_X101Y124_SLICE_X158Y124_CO6),
.I3(CLBLL_L_X102Y126_SLICE_X161Y126_D5Q),
.I4(CLBLM_R_X101Y128_SLICE_X158Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y124_SLICE_X159Y124_AO5),
.O6(CLBLM_R_X101Y124_SLICE_X159Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y125_SLICE_X158Y125_BO5),
.Q(CLBLM_R_X101Y125_SLICE_X158Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y125_SLICE_X158Y125_AO6),
.Q(CLBLM_R_X101Y125_SLICE_X158Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y125_SLICE_X158Y125_BO6),
.Q(CLBLM_R_X101Y125_SLICE_X158Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f1f0f1f5f1f5f1f)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(1'b1),
.I5(CLBLL_L_X100Y125_SLICE_X157Y125_C5Q),
.O5(CLBLM_R_X101Y125_SLICE_X158Y125_DO5),
.O6(CLBLM_R_X101Y125_SLICE_X158Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(CLBLM_R_X101Y125_SLICE_X158Y125_AQ),
.I2(CLBLL_L_X100Y125_SLICE_X157Y125_A5Q),
.I3(CLBLM_R_X101Y125_SLICE_X158Y125_BQ),
.I4(CLBLM_R_X101Y125_SLICE_X158Y125_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y125_SLICE_X158Y125_CO5),
.O6(CLBLM_R_X101Y125_SLICE_X158Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y125_SLICE_X158Y125_BQ),
.I2(CLBLM_R_X101Y125_SLICE_X158Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y125_SLICE_X158Y125_BO5),
.O6(CLBLM_R_X101Y125_SLICE_X158Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4055405551555155)
  ) CLBLM_R_X101Y125_SLICE_X158Y125_ALUT (
.I0(CLBLM_R_X101Y125_SLICE_X158Y125_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y126_SLICE_X158Y126_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(1'b1),
.I5(CLBLM_R_X101Y125_SLICE_X158Y125_CO6),
.O5(CLBLM_R_X101Y125_SLICE_X158Y125_AO5),
.O6(CLBLM_R_X101Y125_SLICE_X158Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y125_SLICE_X159Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y125_SLICE_X159Y125_DO5),
.O6(CLBLM_R_X101Y125_SLICE_X159Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y125_SLICE_X159Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y125_SLICE_X159Y125_CO5),
.O6(CLBLM_R_X101Y125_SLICE_X159Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y125_SLICE_X159Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y125_SLICE_X159Y125_BO5),
.O6(CLBLM_R_X101Y125_SLICE_X159Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y125_SLICE_X159Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y125_SLICE_X159Y125_AO5),
.O6(CLBLM_R_X101Y125_SLICE_X159Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y126_SLICE_X158Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y126_SLICE_X158Y126_AO5),
.Q(CLBLM_R_X101Y126_SLICE_X158Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y126_SLICE_X158Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y126_SLICE_X158Y126_AO6),
.Q(CLBLM_R_X101Y126_SLICE_X158Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y126_SLICE_X158Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X158Y126_DO5),
.O6(CLBLM_R_X101Y126_SLICE_X158Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y126_SLICE_X158Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X158Y126_CO5),
.O6(CLBLM_R_X101Y126_SLICE_X158Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555f5f55557777)
  ) CLBLM_R_X101Y126_SLICE_X158Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X100Y124_SLICE_X157Y124_B5Q),
.I3(1'b1),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y126_SLICE_X158Y126_BO5),
.O6(CLBLM_R_X101Y126_SLICE_X158Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X101Y126_SLICE_X158Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y126_SLICE_X158Y126_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X103Y125_SLICE_X162Y125_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X158Y126_AO5),
.O6(CLBLM_R_X101Y126_SLICE_X158Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y126_SLICE_X159Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y126_SLICE_X159Y126_AO5),
.Q(CLBLM_R_X101Y126_SLICE_X159Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y126_SLICE_X159Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y126_SLICE_X159Y126_AO6),
.Q(CLBLM_R_X101Y126_SLICE_X159Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y126_SLICE_X159Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X159Y126_DO5),
.O6(CLBLM_R_X101Y126_SLICE_X159Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y126_SLICE_X159Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X159Y126_CO5),
.O6(CLBLM_R_X101Y126_SLICE_X159Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y126_SLICE_X159Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X159Y126_BO5),
.O6(CLBLM_R_X101Y126_SLICE_X159Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88228822a0a00a0a)
  ) CLBLM_R_X101Y126_SLICE_X159Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y127_SLICE_X159Y127_A5Q),
.I2(CLBLM_R_X101Y126_SLICE_X159Y126_AQ),
.I3(CLBLM_L_X98Y125_SLICE_X155Y125_A5Q),
.I4(CLBLL_L_X100Y124_SLICE_X156Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y126_SLICE_X159Y126_AO5),
.O6(CLBLM_R_X101Y126_SLICE_X159Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y127_SLICE_X158Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X158Y127_DO5),
.O6(CLBLM_R_X101Y127_SLICE_X158Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y127_SLICE_X158Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X158Y127_CO5),
.O6(CLBLM_R_X101Y127_SLICE_X158Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y127_SLICE_X158Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X158Y127_BO5),
.O6(CLBLM_R_X101Y127_SLICE_X158Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y127_SLICE_X158Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X158Y127_AO5),
.O6(CLBLM_R_X101Y127_SLICE_X158Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y127_SLICE_X159Y127_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y127_SLICE_X159Y127_AO5),
.Q(CLBLM_R_X101Y127_SLICE_X159Y127_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y127_SLICE_X159Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y127_SLICE_X159Y127_AO6),
.Q(CLBLM_R_X101Y127_SLICE_X159Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y127_SLICE_X159Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X159Y127_DO5),
.O6(CLBLM_R_X101Y127_SLICE_X159Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y127_SLICE_X159Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X159Y127_CO5),
.O6(CLBLM_R_X101Y127_SLICE_X159Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2e2d1e2d1d1e2)
  ) CLBLM_R_X101Y127_SLICE_X159Y127_BLUT (
.I0(CLBLL_L_X102Y127_SLICE_X160Y127_CQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y127_SLICE_X159Y127_AQ),
.I3(CLBLL_L_X102Y129_SLICE_X160Y129_CQ),
.I4(CLBLL_L_X102Y127_SLICE_X160Y127_C5Q),
.I5(CLBLL_L_X102Y127_SLICE_X160Y127_BQ),
.O5(CLBLM_R_X101Y127_SLICE_X159Y127_BO5),
.O6(CLBLM_R_X101Y127_SLICE_X159Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88882222a00aa00a)
  ) CLBLM_R_X101Y127_SLICE_X159Y127_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X100Y129_SLICE_X156Y129_AQ),
.I2(CLBLM_R_X101Y127_SLICE_X159Y127_AQ),
.I3(CLBLM_L_X98Y126_SLICE_X155Y126_A5Q),
.I4(CLBLM_R_X97Y126_SLICE_X153Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y127_SLICE_X159Y127_AO5),
.O6(CLBLM_R_X101Y127_SLICE_X159Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y128_SLICE_X158Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y128_SLICE_X158Y128_AO5),
.Q(CLBLM_R_X101Y128_SLICE_X158Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y128_SLICE_X158Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y128_SLICE_X158Y128_AO6),
.Q(CLBLM_R_X101Y128_SLICE_X158Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X158Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X158Y128_DO5),
.O6(CLBLM_R_X101Y128_SLICE_X158Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X158Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X158Y128_CO5),
.O6(CLBLM_R_X101Y128_SLICE_X158Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X158Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X158Y128_BO5),
.O6(CLBLM_R_X101Y128_SLICE_X158Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa82828282)
  ) CLBLM_R_X101Y128_SLICE_X158Y128_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y129_SLICE_X158Y129_B5Q),
.I2(CLBLL_L_X100Y129_SLICE_X157Y129_A5Q),
.I3(1'b1),
.I4(CLBLL_L_X100Y126_SLICE_X157Y126_DO6),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X158Y128_AO5),
.O6(CLBLM_R_X101Y128_SLICE_X158Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X159Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X159Y128_DO5),
.O6(CLBLM_R_X101Y128_SLICE_X159Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X159Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X159Y128_CO5),
.O6(CLBLM_R_X101Y128_SLICE_X159Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X159Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X159Y128_BO5),
.O6(CLBLM_R_X101Y128_SLICE_X159Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y128_SLICE_X159Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y128_SLICE_X159Y128_AO5),
.O6(CLBLM_R_X101Y128_SLICE_X159Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y129_SLICE_X158Y129_AO5),
.Q(CLBLM_R_X101Y129_SLICE_X158Y129_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y129_SLICE_X158Y129_BO5),
.Q(CLBLM_R_X101Y129_SLICE_X158Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y129_SLICE_X158Y129_AO6),
.Q(CLBLM_R_X101Y129_SLICE_X158Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y129_SLICE_X158Y129_BO6),
.Q(CLBLM_R_X101Y129_SLICE_X158Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_DLUT (
.I0(CLBLM_R_X101Y129_SLICE_X159Y129_AQ),
.I1(CLBLM_R_X101Y129_SLICE_X158Y129_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y129_SLICE_X158Y129_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X101Y130_SLICE_X158Y130_C5Q),
.O5(CLBLM_R_X101Y129_SLICE_X158Y129_DO5),
.O6(CLBLM_R_X101Y129_SLICE_X158Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_CLUT (
.I0(CLBLM_R_X101Y129_SLICE_X158Y129_BQ),
.I1(CLBLM_R_X101Y130_SLICE_X158Y130_BQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y130_SLICE_X158Y130_CQ),
.I4(CLBLM_R_X101Y129_SLICE_X158Y129_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y129_SLICE_X158Y129_CO5),
.O6(CLBLM_R_X101Y129_SLICE_X158Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y129_SLICE_X158Y129_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y130_SLICE_X158Y130_CQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y129_SLICE_X158Y129_BO5),
.O6(CLBLM_R_X101Y129_SLICE_X158Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X101Y129_SLICE_X158Y129_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y129_SLICE_X158Y129_AQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y129_SLICE_X159Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y129_SLICE_X158Y129_AO5),
.O6(CLBLM_R_X101Y129_SLICE_X158Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y129_SLICE_X159Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y129_SLICE_X159Y129_AO6),
.Q(CLBLM_R_X101Y129_SLICE_X159Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y129_SLICE_X159Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y129_SLICE_X159Y129_DO5),
.O6(CLBLM_R_X101Y129_SLICE_X159Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y129_SLICE_X159Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y129_SLICE_X159Y129_CO5),
.O6(CLBLM_R_X101Y129_SLICE_X159Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00441155ffffffff)
  ) CLBLM_R_X101Y129_SLICE_X159Y129_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(1'b1),
.I3(CLBLL_L_X100Y129_SLICE_X157Y129_A5Q),
.I4(RIOB33_X105Y137_IOB_X1Y138_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y129_SLICE_X159Y129_BO5),
.O6(CLBLM_R_X101Y129_SLICE_X159Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h008f00bf008f00bf)
  ) CLBLM_R_X101Y129_SLICE_X159Y129_ALUT (
.I0(CLBLL_L_X102Y129_SLICE_X160Y129_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X101Y129_SLICE_X159Y129_BO6),
.I4(CLBLM_R_X101Y129_SLICE_X158Y129_DO6),
.I5(1'b1),
.O5(CLBLM_R_X101Y129_SLICE_X159Y129_AO5),
.O6(CLBLM_R_X101Y129_SLICE_X159Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X158Y130_AO5),
.Q(CLBLM_R_X101Y130_SLICE_X158Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X158Y130_CO5),
.Q(CLBLM_R_X101Y130_SLICE_X158Y130_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X158Y130_AO6),
.Q(CLBLM_R_X101Y130_SLICE_X158Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X158Y130_BO6),
.Q(CLBLM_R_X101Y130_SLICE_X158Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X158Y130_CO6),
.Q(CLBLM_R_X101Y130_SLICE_X158Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h01ff01ff31ff31ff)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_DLUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(CLBLM_R_X101Y128_SLICE_X158Y128_A5Q),
.O5(CLBLM_R_X101Y130_SLICE_X158Y130_DO5),
.O6(CLBLM_R_X101Y130_SLICE_X158Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y129_SLICE_X158Y129_A5Q),
.I2(CLBLM_R_X101Y130_SLICE_X158Y130_BQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y130_SLICE_X158Y130_CO5),
.O6(CLBLM_R_X101Y130_SLICE_X158Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5515051555150515)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_BLUT (
.I0(CLBLM_R_X101Y130_SLICE_X158Y130_DO6),
.I1(CLBLM_R_X101Y129_SLICE_X158Y129_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLL_L_X102Y129_SLICE_X160Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y130_SLICE_X158Y130_BO5),
.O6(CLBLM_R_X101Y130_SLICE_X158Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X101Y130_SLICE_X158Y130_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y130_SLICE_X158Y130_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y130_SLICE_X160Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y130_SLICE_X158Y130_AO5),
.O6(CLBLM_R_X101Y130_SLICE_X158Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X159Y130_BO5),
.Q(CLBLM_R_X101Y130_SLICE_X159Y130_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X159Y130_AO6),
.Q(CLBLM_R_X101Y130_SLICE_X159Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y130_SLICE_X159Y130_BO6),
.Q(CLBLM_R_X101Y130_SLICE_X159Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb8b88bb88b8bb8)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_DLUT (
.I0(CLBLM_L_X98Y131_SLICE_X155Y131_DQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y130_SLICE_X159Y130_BQ),
.I3(CLBLM_R_X101Y130_SLICE_X159Y130_AQ),
.I4(CLBLM_R_X101Y130_SLICE_X159Y130_B5Q),
.I5(CLBLM_R_X101Y131_SLICE_X159Y131_A5Q),
.O5(CLBLM_R_X101Y130_SLICE_X159Y130_DO5),
.O6(CLBLM_R_X101Y130_SLICE_X159Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_CLUT (
.I0(CLBLL_L_X102Y130_SLICE_X160Y130_AQ),
.I1(CLBLM_R_X101Y131_SLICE_X159Y131_A5Q),
.I2(CLBLM_R_X101Y130_SLICE_X159Y130_BQ),
.I3(CLBLM_R_X101Y130_SLICE_X159Y130_AQ),
.I4(CLBLM_R_X101Y130_SLICE_X159Y130_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y130_SLICE_X159Y130_CO5),
.O6(CLBLM_R_X101Y130_SLICE_X159Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y130_SLICE_X159Y130_BQ),
.I2(CLBLM_R_X101Y130_SLICE_X159Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y130_SLICE_X159Y130_BO5),
.O6(CLBLM_R_X101Y130_SLICE_X159Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbea514000000000)
  ) CLBLM_R_X101Y130_SLICE_X159Y130_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y131_SLICE_X159Y131_DQ),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(CLBLM_R_X101Y130_SLICE_X159Y130_CO6),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y130_SLICE_X159Y130_AO5),
.O6(CLBLM_R_X101Y130_SLICE_X159Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X158Y131_BO5),
.Q(CLBLM_R_X101Y131_SLICE_X158Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X158Y131_AO6),
.Q(CLBLM_R_X101Y131_SLICE_X158Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X158Y131_BO6),
.Q(CLBLM_R_X101Y131_SLICE_X158Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_DLUT (
.I0(CLBLM_R_X101Y131_SLICE_X159Y131_AQ),
.I1(CLBLM_R_X101Y131_SLICE_X158Y131_AQ),
.I2(CLBLM_L_X98Y131_SLICE_X155Y131_D5Q),
.I3(CLBLM_R_X101Y131_SLICE_X158Y131_BQ),
.I4(CLBLM_R_X101Y131_SLICE_X158Y131_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y131_SLICE_X158Y131_DO5),
.O6(CLBLM_R_X101Y131_SLICE_X158Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_CLUT (
.I0(CLBLM_R_X101Y131_SLICE_X159Y131_AQ),
.I1(CLBLM_R_X101Y131_SLICE_X158Y131_AQ),
.I2(CLBLM_R_X101Y130_SLICE_X158Y130_A5Q),
.I3(CLBLM_R_X101Y131_SLICE_X158Y131_BQ),
.I4(CLBLM_R_X101Y131_SLICE_X158Y131_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y131_SLICE_X158Y131_CO5),
.O6(CLBLM_R_X101Y131_SLICE_X158Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y131_SLICE_X158Y131_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X101Y131_SLICE_X159Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y131_SLICE_X158Y131_BO5),
.O6(CLBLM_R_X101Y131_SLICE_X158Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d800000000)
  ) CLBLM_R_X101Y131_SLICE_X158Y131_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y131_SLICE_X159Y131_D5Q),
.I2(RIOB33_X105Y125_IOB_X1Y126_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X101Y131_SLICE_X158Y131_CO6),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y131_SLICE_X158Y131_AO5),
.O6(CLBLM_R_X101Y131_SLICE_X158Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_AO5),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_BO5),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_CO5),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_DO5),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_AO6),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_BO6),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_CO6),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y131_SLICE_X159Y131_DO6),
.Q(CLBLM_R_X101Y131_SLICE_X159Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0000cc84848484)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_DLUT (
.I0(CLBLM_R_X101Y131_SLICE_X159Y131_DQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y131_SLICE_X158Y131_B5Q),
.I3(CLBLM_R_X101Y131_SLICE_X159Y131_A5Q),
.I4(CLBLM_R_X101Y131_SLICE_X159Y131_CQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y131_SLICE_X159Y131_DO5),
.O6(CLBLM_R_X101Y131_SLICE_X159Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00cc00c48488484)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_CLUT (
.I0(CLBLM_R_X101Y133_SLICE_X159Y133_AQ),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y128_SLICE_X158Y128_A5Q),
.I3(CLBLL_L_X102Y131_SLICE_X160Y131_B5Q),
.I4(CLBLM_R_X101Y131_SLICE_X159Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y131_SLICE_X159Y131_CO5),
.O6(CLBLM_R_X101Y131_SLICE_X159Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_BLUT (
.I0(CLBLM_R_X101Y132_SLICE_X159Y132_B5Q),
.I1(CLBLL_L_X102Y131_SLICE_X160Y131_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y131_SLICE_X159Y131_BO5),
.O6(CLBLM_R_X101Y131_SLICE_X159Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_R_X101Y131_SLICE_X159Y131_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y130_SLICE_X159Y130_B5Q),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y131_SLICE_X158Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y131_SLICE_X159Y131_AO5),
.O6(CLBLM_R_X101Y131_SLICE_X159Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y132_SLICE_X158Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y132_SLICE_X158Y132_AO5),
.Q(CLBLM_R_X101Y132_SLICE_X158Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y132_SLICE_X158Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y132_SLICE_X158Y132_AO6),
.Q(CLBLM_R_X101Y132_SLICE_X158Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y132_SLICE_X158Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y132_SLICE_X158Y132_DO5),
.O6(CLBLM_R_X101Y132_SLICE_X158Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y132_SLICE_X158Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y132_SLICE_X158Y132_CO5),
.O6(CLBLM_R_X101Y132_SLICE_X158Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y132_SLICE_X158Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y132_SLICE_X158Y132_BO5),
.O6(CLBLM_R_X101Y132_SLICE_X158Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X101Y132_SLICE_X158Y132_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y132_SLICE_X158Y132_A5Q),
.I2(CLBLM_R_X101Y130_SLICE_X158Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y132_SLICE_X158Y132_AO5),
.O6(CLBLM_R_X101Y132_SLICE_X158Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y132_SLICE_X159Y132_BO5),
.Q(CLBLM_R_X101Y132_SLICE_X159Y132_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y132_SLICE_X159Y132_AO6),
.Q(CLBLM_R_X101Y132_SLICE_X159Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y132_SLICE_X159Y132_BO6),
.Q(CLBLM_R_X101Y132_SLICE_X159Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_DLUT (
.I0(CLBLM_L_X98Y130_SLICE_X155Y130_D5Q),
.I1(CLBLM_R_X101Y131_SLICE_X159Y131_B5Q),
.I2(CLBLM_R_X101Y132_SLICE_X159Y132_BQ),
.I3(CLBLM_R_X101Y132_SLICE_X159Y132_AQ),
.I4(CLBLM_R_X101Y132_SLICE_X159Y132_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y132_SLICE_X159Y132_DO5),
.O6(CLBLM_R_X101Y132_SLICE_X159Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeebebbe14414114)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y131_SLICE_X159Y131_B5Q),
.I2(CLBLM_R_X101Y132_SLICE_X159Y132_BQ),
.I3(CLBLM_R_X101Y132_SLICE_X159Y132_AQ),
.I4(CLBLM_R_X101Y132_SLICE_X159Y132_B5Q),
.I5(CLBLM_R_X101Y132_SLICE_X158Y132_A5Q),
.O5(CLBLM_R_X101Y132_SLICE_X159Y132_CO5),
.O6(CLBLM_R_X101Y132_SLICE_X159Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y132_SLICE_X159Y132_BQ),
.I2(CLBLM_R_X101Y132_SLICE_X159Y132_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y132_SLICE_X159Y132_BO5),
.O6(CLBLM_R_X101Y132_SLICE_X159Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbea514000000000)
  ) CLBLM_R_X101Y132_SLICE_X159Y132_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y131_SLICE_X159Y131_C5Q),
.I3(RIOB33_X105Y139_IOB_X1Y140_I),
.I4(CLBLM_R_X101Y132_SLICE_X159Y132_CO6),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y132_SLICE_X159Y132_AO5),
.O6(CLBLM_R_X101Y132_SLICE_X159Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y133_SLICE_X158Y133_BO5),
.Q(CLBLM_R_X101Y133_SLICE_X158Y133_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y133_SLICE_X158Y133_AO6),
.Q(CLBLM_R_X101Y133_SLICE_X158Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y133_SLICE_X158Y133_BO6),
.Q(CLBLM_R_X101Y133_SLICE_X158Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3cc3c33c)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_DLUT (
.I0(CLBLM_L_X98Y132_SLICE_X155Y132_CQ),
.I1(CLBLM_R_X101Y133_SLICE_X158Y133_AQ),
.I2(CLBLM_R_X101Y134_SLICE_X158Y134_A5Q),
.I3(CLBLM_R_X101Y133_SLICE_X158Y133_BQ),
.I4(CLBLM_R_X101Y133_SLICE_X158Y133_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X101Y133_SLICE_X158Y133_DO5),
.O6(CLBLM_R_X101Y133_SLICE_X158Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caac3aac3aa3c)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_CLUT (
.I0(CLBLM_R_X101Y130_SLICE_X158Y130_AQ),
.I1(CLBLM_R_X101Y133_SLICE_X158Y133_AQ),
.I2(CLBLM_R_X101Y133_SLICE_X158Y133_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X101Y133_SLICE_X158Y133_B5Q),
.I5(CLBLM_R_X101Y134_SLICE_X158Y134_A5Q),
.O5(CLBLM_R_X101Y133_SLICE_X158Y133_CO5),
.O6(CLBLM_R_X101Y133_SLICE_X158Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X101Y133_SLICE_X158Y133_BQ),
.I2(CLBLM_R_X101Y133_SLICE_X158Y133_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y133_SLICE_X158Y133_BO5),
.O6(CLBLM_R_X101Y133_SLICE_X158Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa8aa2000a80020)
  ) CLBLM_R_X101Y133_SLICE_X158Y133_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X101Y133_SLICE_X159Y133_AQ),
.I5(CLBLM_R_X101Y133_SLICE_X158Y133_CO6),
.O5(CLBLM_R_X101Y133_SLICE_X158Y133_AO5),
.O6(CLBLM_R_X101Y133_SLICE_X158Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y133_SLICE_X159Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y133_SLICE_X159Y133_AO5),
.Q(CLBLM_R_X101Y133_SLICE_X159Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y133_SLICE_X159Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y133_SLICE_X159Y133_AO6),
.Q(CLBLM_R_X101Y133_SLICE_X159Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y133_SLICE_X159Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y133_SLICE_X159Y133_DO5),
.O6(CLBLM_R_X101Y133_SLICE_X159Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y133_SLICE_X159Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y133_SLICE_X159Y133_CO5),
.O6(CLBLM_R_X101Y133_SLICE_X159Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f909f909f606)
  ) CLBLM_R_X101Y133_SLICE_X159Y133_BLUT (
.I0(CLBLM_R_X101Y135_SLICE_X159Y135_A5Q),
.I1(CLBLM_R_X101Y134_SLICE_X159Y134_CQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLL_L_X100Y133_SLICE_X156Y133_AQ),
.I4(CLBLM_R_X101Y134_SLICE_X159Y134_AQ),
.I5(CLBLM_R_X101Y134_SLICE_X159Y134_C5Q),
.O5(CLBLM_R_X101Y133_SLICE_X159Y133_BO5),
.O6(CLBLM_R_X101Y133_SLICE_X159Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc030c030a0a05050)
  ) CLBLM_R_X101Y133_SLICE_X159Y133_ALUT (
.I0(CLBLL_L_X100Y134_SLICE_X156Y134_A5Q),
.I1(CLBLM_R_X101Y134_SLICE_X158Y134_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X101Y131_SLICE_X159Y131_D5Q),
.I4(CLBLM_R_X101Y131_SLICE_X159Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y133_SLICE_X159Y133_AO5),
.O6(CLBLM_R_X101Y133_SLICE_X159Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y134_SLICE_X158Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y134_SLICE_X158Y134_AO5),
.Q(CLBLM_R_X101Y134_SLICE_X158Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y134_SLICE_X158Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y134_SLICE_X158Y134_AO6),
.Q(CLBLM_R_X101Y134_SLICE_X158Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y134_SLICE_X158Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y134_SLICE_X158Y134_DO5),
.O6(CLBLM_R_X101Y134_SLICE_X158Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y134_SLICE_X158Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y134_SLICE_X158Y134_CO5),
.O6(CLBLM_R_X101Y134_SLICE_X158Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed1221edde2112)
  ) CLBLM_R_X101Y134_SLICE_X158Y134_BLUT (
.I0(CLBLL_L_X100Y134_SLICE_X156Y134_A5Q),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y134_SLICE_X158Y134_AQ),
.I3(CLBLM_R_X101Y134_SLICE_X159Y134_BQ),
.I4(CLBLM_R_X101Y132_SLICE_X158Y132_AQ),
.I5(CLBLL_L_X100Y134_SLICE_X156Y134_AQ),
.O5(CLBLM_R_X101Y134_SLICE_X158Y134_BO5),
.O6(CLBLM_R_X101Y134_SLICE_X158Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_R_X101Y134_SLICE_X158Y134_ALUT (
.I0(CLBLM_R_X101Y133_SLICE_X158Y133_B5Q),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X101Y134_SLICE_X159Y134_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y134_SLICE_X158Y134_AO5),
.O6(CLBLM_R_X101Y134_SLICE_X158Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y134_SLICE_X159Y134_CO5),
.Q(CLBLM_R_X101Y134_SLICE_X159Y134_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y134_SLICE_X159Y134_AO6),
.Q(CLBLM_R_X101Y134_SLICE_X159Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y134_SLICE_X159Y134_BO6),
.Q(CLBLM_R_X101Y134_SLICE_X159Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y134_SLICE_X159Y134_CO6),
.Q(CLBLM_R_X101Y134_SLICE_X159Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff699600006996)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_DLUT (
.I0(CLBLM_R_X101Y134_SLICE_X159Y134_C5Q),
.I1(CLBLM_R_X101Y134_SLICE_X159Y134_CQ),
.I2(CLBLM_R_X101Y135_SLICE_X159Y135_A5Q),
.I3(CLBLM_R_X101Y134_SLICE_X159Y134_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLL_L_X102Y134_SLICE_X160Y134_A5Q),
.O5(CLBLM_R_X101Y134_SLICE_X159Y134_DO5),
.O6(CLBLM_R_X101Y134_SLICE_X159Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y134_SLICE_X159Y134_CQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y134_SLICE_X159Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y134_SLICE_X159Y134_CO5),
.O6(CLBLM_R_X101Y134_SLICE_X159Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc5000000000)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y134_SLICE_X158Y134_BO6),
.I2(RIOB33_X105Y141_IOB_X1Y141_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X101Y133_SLICE_X159Y133_A5Q),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y134_SLICE_X159Y134_BO5),
.O6(CLBLM_R_X101Y134_SLICE_X159Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3c000000000)
  ) CLBLM_R_X101Y134_SLICE_X159Y134_ALUT (
.I0(CLBLM_R_X101Y134_SLICE_X159Y134_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y135_SLICE_X159Y135_DQ),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X101Y134_SLICE_X159Y134_AO5),
.O6(CLBLM_R_X101Y134_SLICE_X159Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X158Y135_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X158Y135_AO5),
.Q(CLBLM_R_X101Y135_SLICE_X158Y135_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X158Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X158Y135_AO6),
.Q(CLBLM_R_X101Y135_SLICE_X158Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y135_SLICE_X158Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X158Y135_DO5),
.O6(CLBLM_R_X101Y135_SLICE_X158Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y135_SLICE_X158Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X158Y135_CO5),
.O6(CLBLM_R_X101Y135_SLICE_X158Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14eb41eb41be14)
  ) CLBLM_R_X101Y135_SLICE_X158Y135_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X102Y135_SLICE_X160Y135_AQ),
.I2(CLBLM_R_X101Y135_SLICE_X158Y135_AQ),
.I3(CLBLL_L_X100Y133_SLICE_X156Y133_A5Q),
.I4(CLBLM_R_X101Y135_SLICE_X159Y135_AQ),
.I5(CLBLM_R_X101Y135_SLICE_X158Y135_A5Q),
.O5(CLBLM_R_X101Y135_SLICE_X158Y135_BO5),
.O6(CLBLM_R_X101Y135_SLICE_X158Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X101Y135_SLICE_X158Y135_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y135_SLICE_X158Y135_AQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y135_SLICE_X159Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X158Y135_AO5),
.O6(CLBLM_R_X101Y135_SLICE_X158Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_AO5),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_BO5),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_CO5),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_DO5),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_AO6),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_BO6),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_CO6),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y135_SLICE_X159Y135_DO6),
.Q(CLBLM_R_X101Y135_SLICE_X159Y135_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa005500c300c300)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_DLUT (
.I0(CLBLM_R_X101Y135_SLICE_X159Y135_C5Q),
.I1(CLBLM_R_X101Y135_SLICE_X158Y135_A5Q),
.I2(CLBLM_R_X101Y135_SLICE_X159Y135_DQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y135_SLICE_X159Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X159Y135_DO5),
.O6(CLBLM_R_X101Y135_SLICE_X159Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa005500c300c300)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_CLUT (
.I0(CLBLM_R_X101Y133_SLICE_X159Y133_A5Q),
.I1(CLBLM_R_X101Y135_SLICE_X159Y135_CQ),
.I2(CLBLL_L_X102Y136_SLICE_X160Y136_B5Q),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X101Y135_SLICE_X159Y135_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X159Y135_CO5),
.O6(CLBLM_R_X101Y135_SLICE_X159Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y136_SLICE_X159Y136_B5Q),
.I3(1'b1),
.I4(CLBLL_L_X102Y136_SLICE_X160Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X159Y135_BO5),
.O6(CLBLM_R_X101Y135_SLICE_X159Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X101Y135_SLICE_X159Y135_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X101Y134_SLICE_X159Y134_C5Q),
.I3(CLBLL_L_X102Y135_SLICE_X160Y135_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y135_SLICE_X159Y135_AO5),
.O6(CLBLM_R_X101Y135_SLICE_X159Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y136_SLICE_X158Y136_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y136_SLICE_X158Y136_AO5),
.Q(CLBLM_R_X101Y136_SLICE_X158Y136_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y136_SLICE_X158Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y136_SLICE_X158Y136_AO6),
.Q(CLBLM_R_X101Y136_SLICE_X158Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y136_SLICE_X158Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y136_SLICE_X158Y136_DO5),
.O6(CLBLM_R_X101Y136_SLICE_X158Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y136_SLICE_X158Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y136_SLICE_X158Y136_CO5),
.O6(CLBLM_R_X101Y136_SLICE_X158Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y136_SLICE_X158Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y136_SLICE_X158Y136_BO5),
.O6(CLBLM_R_X101Y136_SLICE_X158Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X101Y136_SLICE_X158Y136_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X101Y132_SLICE_X158Y132_AQ),
.I3(1'b1),
.I4(CLBLM_R_X101Y136_SLICE_X158Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X101Y136_SLICE_X158Y136_AO5),
.O6(CLBLM_R_X101Y136_SLICE_X158Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y136_SLICE_X159Y136_BO5),
.Q(CLBLM_R_X101Y136_SLICE_X159Y136_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y136_SLICE_X159Y136_AO6),
.Q(CLBLM_R_X101Y136_SLICE_X159Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X101Y136_SLICE_X159Y136_BO6),
.Q(CLBLM_R_X101Y136_SLICE_X159Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb8b88bb88b8bb8)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_DLUT (
.I0(CLBLL_L_X100Y134_SLICE_X156Y134_BQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X101Y135_SLICE_X159Y135_B5Q),
.I3(CLBLM_R_X101Y136_SLICE_X159Y136_BQ),
.I4(CLBLM_R_X101Y136_SLICE_X159Y136_B5Q),
.I5(CLBLM_R_X101Y136_SLICE_X159Y136_AQ),
.O5(CLBLM_R_X101Y136_SLICE_X159Y136_DO5),
.O6(CLBLM_R_X101Y136_SLICE_X159Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd8d88dd88d8dd8)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X101Y136_SLICE_X158Y136_A5Q),
.I2(CLBLM_R_X101Y135_SLICE_X159Y135_B5Q),
.I3(CLBLM_R_X101Y136_SLICE_X159Y136_BQ),
.I4(CLBLM_R_X101Y136_SLICE_X159Y136_B5Q),
.I5(CLBLM_R_X101Y136_SLICE_X159Y136_AQ),
.O5(CLBLM_R_X101Y136_SLICE_X159Y136_CO5),
.O6(CLBLM_R_X101Y136_SLICE_X159Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X101Y136_SLICE_X159Y136_BQ),
.I2(CLBLM_R_X101Y136_SLICE_X159Y136_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y136_SLICE_X159Y136_BO5),
.O6(CLBLM_R_X101Y136_SLICE_X159Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e0d0c030201000)
  ) CLBLM_R_X101Y136_SLICE_X159Y136_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X101Y135_SLICE_X159Y135_CQ),
.I5(CLBLM_R_X101Y136_SLICE_X159Y136_CO6),
.O5(CLBLM_R_X101Y136_SLICE_X159Y136_AO5),
.O6(CLBLM_R_X101Y136_SLICE_X159Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_BO5),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_AO5),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_BO6),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_DO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_CLUT (
.I0(CLBLM_R_X103Y112_SLICE_X162Y112_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X103Y111_SLICE_X162Y111_BQ),
.I4(CLBLM_R_X103Y111_SLICE_X162Y111_B5Q),
.I5(CLBLM_R_X101Y111_SLICE_X159Y111_BQ),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_CO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X101Y111_SLICE_X159Y111_BQ),
.I4(CLBLM_R_X103Y111_SLICE_X162Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_BO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05f5fc0c0c0c0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X103Y111_SLICE_X162Y111_AQ),
.I3(1'b1),
.I4(CLBLM_R_X103Y111_SLICE_X162Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_AO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_DO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_CO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_BO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_AO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_BO5),
.Q(CLBLM_R_X103Y112_SLICE_X162Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_CO5),
.Q(CLBLM_R_X103Y112_SLICE_X162Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_BO6),
.Q(CLBLM_R_X103Y112_SLICE_X162Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_CO6),
.Q(CLBLM_R_X103Y112_SLICE_X162Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966969969669)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_DLUT (
.I0(CLBLM_R_X103Y112_SLICE_X162Y112_BQ),
.I1(CLBLM_R_X103Y112_SLICE_X162Y112_CQ),
.I2(CLBLM_R_X101Y111_SLICE_X159Y111_AQ),
.I3(CLBLM_R_X103Y112_SLICE_X162Y112_C5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_DO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_CLUT (
.I0(CLBLM_R_X103Y112_SLICE_X162Y112_BQ),
.I1(CLBLM_R_X103Y112_SLICE_X162Y112_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_CO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cc00cc00)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X103Y111_SLICE_X162Y111_B5Q),
.I4(CLBLM_R_X101Y111_SLICE_X159Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_BO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa555555cc00cc00)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_ALUT (
.I0(CLBLM_R_X103Y112_SLICE_X163Y112_BO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLM_R_X103Y112_SLICE_X163Y112_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_AO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X163Y112_AO5),
.Q(CLBLM_R_X103Y112_SLICE_X163Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y112_SLICE_X163Y112_AO6),
.Q(CLBLM_R_X103Y112_SLICE_X163Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y113_SLICE_X163Y113_BO5),
.Q(CLBLM_R_X103Y112_SLICE_X163Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_DO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_CO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y148_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y112_SLICE_X163Y112_AQ),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_AQ),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_AQ),
.I5(CLBLM_R_X103Y112_SLICE_X163Y112_A5Q),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_BO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X103Y112_SLICE_X163Y112_AQ),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_AO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_AO5),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_BO5),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_AO6),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_BO6),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_DO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55aa55a5aa5)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_CLUT (
.I0(CLBLM_R_X103Y113_SLICE_X162Y113_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q),
.I5(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_CO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_BO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_ALUT (
.I0(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q),
.I1(CLBLL_L_X102Y112_SLICE_X161Y112_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_AO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.Q(CLBLM_R_X103Y113_SLICE_X163Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y114_SLICE_X160Y114_AO5),
.Q(CLBLM_R_X103Y113_SLICE_X163Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_DO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_CO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05fc0c0c0c0)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X103Y113_SLICE_X163Y113_AQ),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_BO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5500ffcccc0000)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(1'b1),
.I3(CLBLL_L_X102Y114_SLICE_X161Y114_BO6),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y116_SLICE_X162Y116_BO5),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y116_SLICE_X162Y116_AO6),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y116_SLICE_X162Y116_BO6),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I2(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X103Y116_SLICE_X162Y116_B5Q),
.I5(CLBLL_L_X102Y117_SLICE_X161Y117_D5Q),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_DO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c639c63939c6)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I2(CLBLL_L_X102Y117_SLICE_X161Y117_B5Q),
.I3(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.I4(CLBLM_R_X103Y116_SLICE_X162Y116_B5Q),
.I5(CLBLL_L_X102Y117_SLICE_X161Y117_D5Q),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_CO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.I2(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_BO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a8080aa0aa000)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y117_SLICE_X161Y117_B5Q),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X103Y116_SLICE_X162Y116_DO6),
.I4(CLBLM_R_X97Y118_SLICE_X153Y118_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_AO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_DO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_CO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_BO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_AO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y117_SLICE_X162Y117_BO5),
.Q(CLBLM_R_X103Y117_SLICE_X162Y117_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y117_SLICE_X162Y117_AO6),
.Q(CLBLM_R_X103Y117_SLICE_X162Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y117_SLICE_X162Y117_BO6),
.Q(CLBLM_R_X103Y117_SLICE_X162Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y117_SLICE_X162Y117_AQ),
.I2(CLBLM_R_X103Y117_SLICE_X162Y117_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X103Y117_SLICE_X162Y117_B5Q),
.I5(CLBLL_L_X102Y117_SLICE_X161Y117_DQ),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_DO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c9c639c63639c)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_CLUT (
.I0(CLBLL_L_X102Y117_SLICE_X161Y117_BQ),
.I1(CLBLM_R_X103Y117_SLICE_X162Y117_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X103Y117_SLICE_X162Y117_BQ),
.I4(CLBLM_R_X103Y117_SLICE_X162Y117_B5Q),
.I5(CLBLL_L_X102Y117_SLICE_X161Y117_DQ),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_CO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y117_SLICE_X162Y117_BQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y117_SLICE_X161Y117_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_BO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8aa08aaa8000800)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y117_SLICE_X162Y117_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLL_L_X102Y117_SLICE_X161Y117_BQ),
.I5(CLBLM_R_X97Y118_SLICE_X152Y118_DO6),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_AO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_DO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_CO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_BO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_AO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLL_L_X102Y118_SLICE_X160Y118_AO5),
.Q(CLBLM_R_X103Y119_SLICE_X162Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_DO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_CO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_BO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_AO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y119_SLICE_X163Y119_BO5),
.Q(CLBLM_R_X103Y119_SLICE_X163Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y119_SLICE_X163Y119_AO6),
.Q(CLBLM_R_X103Y119_SLICE_X163Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y119_SLICE_X163Y119_BO6),
.Q(CLBLM_R_X103Y119_SLICE_X163Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y119_SLICE_X163Y119_BQ),
.I3(CLBLM_R_X103Y119_SLICE_X163Y119_AQ),
.I4(CLBLM_R_X103Y119_SLICE_X163Y119_B5Q),
.I5(CLBLM_R_X103Y120_SLICE_X163Y120_BQ),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_DO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_CLUT (
.I0(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y119_SLICE_X163Y119_BQ),
.I3(CLBLM_R_X103Y119_SLICE_X163Y119_AQ),
.I4(CLBLM_R_X103Y119_SLICE_X163Y119_B5Q),
.I5(CLBLM_R_X103Y120_SLICE_X163Y120_BQ),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_CO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y119_SLICE_X163Y119_BQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y120_SLICE_X163Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_BO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa22a2288800800)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X103Y119_SLICE_X163Y119_DO6),
.I4(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.I5(CLBLL_L_X100Y119_SLICE_X157Y119_DO6),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_AO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X162Y120_AO5),
.Q(CLBLM_R_X103Y120_SLICE_X162Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X162Y120_BO5),
.Q(CLBLM_R_X103Y120_SLICE_X162Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X162Y120_CO5),
.Q(CLBLM_R_X103Y120_SLICE_X162Y120_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X162Y120_AO6),
.Q(CLBLM_R_X103Y120_SLICE_X162Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X162Y120_BO6),
.Q(CLBLM_R_X103Y120_SLICE_X162Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X162Y120_CO6),
.Q(CLBLM_R_X103Y120_SLICE_X162Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y120_SLICE_X162Y120_DO5),
.O6(CLBLM_R_X103Y120_SLICE_X162Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f0f00000)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_CLUT (
.I0(CLBLM_R_X103Y120_SLICE_X162Y120_C5Q),
.I1(1'b1),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y120_SLICE_X162Y120_CO5),
.O6(CLBLM_R_X103Y120_SLICE_X162Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y120_SLICE_X162Y120_CQ),
.I3(CLBLM_R_X103Y120_SLICE_X162Y120_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y120_SLICE_X162Y120_BO5),
.O6(CLBLM_R_X103Y120_SLICE_X162Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X103Y120_SLICE_X162Y120_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y120_SLICE_X162Y120_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X103Y120_SLICE_X162Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y120_SLICE_X162Y120_AO5),
.O6(CLBLM_R_X103Y120_SLICE_X162Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X163Y120_BO5),
.Q(CLBLM_R_X103Y120_SLICE_X163Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X163Y120_AO6),
.Q(CLBLM_R_X103Y120_SLICE_X163Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y120_SLICE_X163Y120_BO6),
.Q(CLBLM_R_X103Y120_SLICE_X163Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699696696996)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_DLUT (
.I0(CLBLM_R_X103Y121_SLICE_X163Y121_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y121_SLICE_X163Y121_A5Q),
.I3(CLBLM_R_X103Y120_SLICE_X163Y120_AQ),
.I4(CLBLM_R_X103Y120_SLICE_X163Y120_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y120_SLICE_X163Y120_DO5),
.O6(CLBLM_R_X103Y120_SLICE_X163Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5a55a96696996)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_CLUT (
.I0(CLBLM_R_X103Y121_SLICE_X163Y121_AQ),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X103Y121_SLICE_X163Y121_A5Q),
.I3(CLBLM_R_X103Y120_SLICE_X163Y120_AQ),
.I4(CLBLM_R_X103Y120_SLICE_X163Y120_B5Q),
.I5(CLBLM_R_X103Y120_SLICE_X162Y120_BQ),
.O5(CLBLM_R_X103Y120_SLICE_X163Y120_CO5),
.O6(CLBLM_R_X103Y120_SLICE_X163Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y119_SLICE_X163Y119_AQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y121_SLICE_X163Y121_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y120_SLICE_X163Y120_BO5),
.O6(CLBLM_R_X103Y120_SLICE_X163Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000c0c0a0a0c0c0)
  ) CLBLM_R_X103Y120_SLICE_X163Y120_ALUT (
.I0(CLBLM_R_X103Y120_SLICE_X163Y120_DO6),
.I1(CLBLL_L_X100Y120_SLICE_X157Y120_CO6),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X103Y120_SLICE_X162Y120_BQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y120_SLICE_X163Y120_AO5),
.O6(CLBLM_R_X103Y120_SLICE_X163Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X162Y121_BO5),
.Q(CLBLM_R_X103Y121_SLICE_X162Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X162Y121_AO6),
.Q(CLBLM_R_X103Y121_SLICE_X162Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X162Y121_BO6),
.Q(CLBLM_R_X103Y121_SLICE_X162Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699696696996)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_DLUT (
.I0(CLBLM_R_X103Y121_SLICE_X162Y121_BQ),
.I1(CLBLM_R_X103Y121_SLICE_X162Y121_AQ),
.I2(CLBLL_L_X102Y121_SLICE_X161Y121_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X103Y121_SLICE_X162Y121_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y121_SLICE_X162Y121_DO5),
.O6(CLBLM_R_X103Y121_SLICE_X162Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696696996)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_CLUT (
.I0(CLBLM_R_X103Y121_SLICE_X162Y121_BQ),
.I1(CLBLM_R_X103Y121_SLICE_X162Y121_AQ),
.I2(CLBLL_L_X102Y121_SLICE_X161Y121_A5Q),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X103Y121_SLICE_X162Y121_B5Q),
.I5(CLBLM_R_X103Y120_SLICE_X162Y120_B5Q),
.O5(CLBLM_R_X103Y121_SLICE_X162Y121_CO5),
.O6(CLBLM_R_X103Y121_SLICE_X162Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y121_SLICE_X162Y121_BQ),
.I2(CLBLM_R_X103Y121_SLICE_X162Y121_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y121_SLICE_X162Y121_BO5),
.O6(CLBLM_R_X103Y121_SLICE_X162Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha808aaaaa8080000)
  ) CLBLM_R_X103Y121_SLICE_X162Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y121_SLICE_X162Y121_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(CLBLM_R_X103Y120_SLICE_X162Y120_B5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLL_L_X100Y121_SLICE_X157Y121_DO6),
.O5(CLBLM_R_X103Y121_SLICE_X162Y121_AO5),
.O6(CLBLM_R_X103Y121_SLICE_X162Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X163Y121_AO5),
.Q(CLBLM_R_X103Y121_SLICE_X163Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X163Y121_BO5),
.Q(CLBLM_R_X103Y121_SLICE_X163Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X163Y121_CO5),
.Q(CLBLM_R_X103Y121_SLICE_X163Y121_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X163Y121_AO6),
.Q(CLBLM_R_X103Y121_SLICE_X163Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X163Y121_BO6),
.Q(CLBLM_R_X103Y121_SLICE_X163Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y121_SLICE_X163Y121_CO6),
.Q(CLBLM_R_X103Y121_SLICE_X163Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696966969)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_DLUT (
.I0(CLBLM_R_X103Y121_SLICE_X163Y121_C5Q),
.I1(CLBLM_R_X103Y121_SLICE_X163Y121_CQ),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_CQ),
.I3(1'b1),
.I4(CLBLM_R_X103Y121_SLICE_X163Y121_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X103Y121_SLICE_X163Y121_DO5),
.O6(CLBLM_R_X103Y121_SLICE_X163Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y121_SLICE_X163Y121_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y121_SLICE_X163Y121_CO5),
.O6(CLBLM_R_X103Y121_SLICE_X163Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaaa0000)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y122_SLICE_X163Y122_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X103Y121_SLICE_X163Y121_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y121_SLICE_X163Y121_BO5),
.O6(CLBLM_R_X103Y121_SLICE_X163Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X103Y121_SLICE_X163Y121_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y121_SLICE_X163Y121_AQ),
.I3(1'b1),
.I4(CLBLM_R_X103Y120_SLICE_X163Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y121_SLICE_X163Y121_AO5),
.O6(CLBLM_R_X103Y121_SLICE_X163Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X162Y122_AO5),
.Q(CLBLM_R_X103Y122_SLICE_X162Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X162Y122_BO5),
.Q(CLBLM_R_X103Y122_SLICE_X162Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X162Y122_AO6),
.Q(CLBLM_R_X103Y122_SLICE_X162Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X162Y122_BO6),
.Q(CLBLM_R_X103Y122_SLICE_X162Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cc33c3cc3)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(CLBLM_R_X103Y122_SLICE_X162Y122_BQ),
.I3(CLBLM_R_X103Y122_SLICE_X162Y122_A5Q),
.I4(CLBLM_R_X103Y122_SLICE_X162Y122_B5Q),
.I5(CLBLM_R_X103Y123_SLICE_X162Y123_BQ),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7750225077fa22fa)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X100Y122_SLICE_X157Y122_C5Q),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X103Y121_SLICE_X163Y121_DO6),
.I5(CLBLL_L_X102Y121_SLICE_X161Y121_CQ),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y122_SLICE_X162Y122_BQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y123_SLICE_X162Y123_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y122_SLICE_X162Y122_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X103Y123_SLICE_X163Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_CO5),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_AO6),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_BO6),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_CO6),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_DLUT (
.I0(CLBLM_R_X103Y122_SLICE_X162Y122_AQ),
.I1(CLBLM_R_X103Y123_SLICE_X163Y123_AQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_A5Q),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_R_X103Y122_SLICE_X163Y122_AQ),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f090909090)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_CLUT (
.I0(CLBLL_L_X102Y122_SLICE_X161Y122_C5Q),
.I1(CLBLM_R_X103Y122_SLICE_X162Y122_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(CLBLM_R_X103Y122_SLICE_X162Y122_CO6),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa88882222)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y122_SLICE_X163Y122_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X102Y121_SLICE_X160Y121_CO6),
.I4(CLBLM_R_X103Y122_SLICE_X163Y122_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000a0a0a0a0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_AQ),
.I3(1'b1),
.I4(CLBLM_R_X103Y122_SLICE_X162Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y123_SLICE_X162Y123_AO5),
.Q(CLBLM_R_X103Y123_SLICE_X162Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y123_SLICE_X162Y123_AO6),
.Q(CLBLM_R_X103Y123_SLICE_X162Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y123_SLICE_X162Y123_BO6),
.Q(CLBLM_R_X103Y123_SLICE_X162Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y123_SLICE_X162Y123_CO6),
.Q(CLBLM_R_X103Y123_SLICE_X162Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_DO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2233223303330333)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_CLUT (
.I0(CLBLM_R_X101Y123_SLICE_X159Y123_AQ),
.I1(CLBLM_R_X103Y123_SLICE_X163Y123_CO6),
.I2(CLBLL_L_X102Y122_SLICE_X161Y122_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_CO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2233003333331133)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_BLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X103Y123_SLICE_X163Y123_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X103Y123_SLICE_X162Y123_A5Q),
.I5(CLBLM_R_X103Y122_SLICE_X162Y122_DO6),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_BO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y123_SLICE_X162Y123_A5Q),
.I2(CLBLM_R_X101Y123_SLICE_X159Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_AO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y123_SLICE_X163Y123_AO6),
.Q(CLBLM_R_X103Y123_SLICE_X163Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_DO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f1f1f1f0f0f3f3f)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_CLUT (
.I0(CLBLL_L_X102Y122_SLICE_X161Y122_C5Q),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(1'b1),
.I4(RIOB33_X105Y125_IOB_X1Y125_I),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_CO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555555555757dfdf)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(1'b1),
.I4(CLBLM_R_X103Y122_SLICE_X163Y122_C5Q),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_BO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0300030f0f0f0f)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y122_SLICE_X163Y122_DO6),
.I2(CLBLM_R_X103Y126_SLICE_X163Y126_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X103Y123_SLICE_X162Y123_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_AO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y124_SLICE_X162Y124_BO5),
.Q(CLBLM_R_X103Y124_SLICE_X162Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y124_SLICE_X162Y124_AO6),
.Q(CLBLM_R_X103Y124_SLICE_X162Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y124_SLICE_X162Y124_BO6),
.Q(CLBLM_R_X103Y124_SLICE_X162Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y124_SLICE_X162Y124_AQ),
.I2(CLBLL_L_X102Y124_SLICE_X161Y124_A5Q),
.I3(CLBLM_R_X103Y124_SLICE_X162Y124_BQ),
.I4(CLBLM_R_X103Y124_SLICE_X162Y124_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y124_SLICE_X162Y124_DO5),
.O6(CLBLM_R_X103Y124_SLICE_X162Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c96c396c3693c)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_CLUT (
.I0(CLBLM_R_X103Y120_SLICE_X162Y120_AQ),
.I1(CLBLM_R_X103Y124_SLICE_X162Y124_AQ),
.I2(CLBLM_R_X103Y124_SLICE_X162Y124_BQ),
.I3(RIOB33_X105Y147_IOB_X1Y147_I),
.I4(CLBLM_R_X103Y124_SLICE_X162Y124_B5Q),
.I5(CLBLL_L_X102Y124_SLICE_X161Y124_A5Q),
.O5(CLBLM_R_X103Y124_SLICE_X162Y124_CO5),
.O6(CLBLM_R_X103Y124_SLICE_X162Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y124_SLICE_X162Y124_BQ),
.I2(CLBLM_R_X103Y124_SLICE_X162Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y124_SLICE_X162Y124_BO5),
.O6(CLBLM_R_X103Y124_SLICE_X162Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a80808a808a808)
  ) CLBLM_R_X103Y124_SLICE_X162Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_L_X98Y123_SLICE_X155Y123_DO6),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X103Y124_SLICE_X162Y124_DO6),
.I4(CLBLM_R_X103Y120_SLICE_X162Y120_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y124_SLICE_X162Y124_AO5),
.O6(CLBLM_R_X103Y124_SLICE_X162Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y124_SLICE_X163Y124_BO5),
.Q(CLBLM_R_X103Y124_SLICE_X163Y124_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y124_SLICE_X163Y124_AO6),
.Q(CLBLM_R_X103Y124_SLICE_X163Y124_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y124_SLICE_X163Y124_BO6),
.Q(CLBLM_R_X103Y124_SLICE_X163Y124_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y124_SLICE_X163Y124_AQ),
.I2(CLBLL_L_X102Y124_SLICE_X160Y124_C5Q),
.I3(CLBLM_R_X103Y124_SLICE_X163Y124_BQ),
.I4(CLBLM_R_X103Y124_SLICE_X163Y124_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y124_SLICE_X163Y124_DO5),
.O6(CLBLM_R_X103Y124_SLICE_X163Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22dd22d2dd2)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLL_L_X102Y124_SLICE_X160Y124_AQ),
.I2(CLBLL_L_X102Y124_SLICE_X160Y124_C5Q),
.I3(CLBLM_R_X103Y124_SLICE_X163Y124_BQ),
.I4(CLBLM_R_X103Y124_SLICE_X163Y124_B5Q),
.I5(CLBLM_R_X103Y124_SLICE_X163Y124_AQ),
.O5(CLBLM_R_X103Y124_SLICE_X163Y124_CO5),
.O6(CLBLM_R_X103Y124_SLICE_X163Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y124_SLICE_X163Y124_BQ),
.I2(CLBLM_R_X103Y124_SLICE_X163Y124_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y124_SLICE_X163Y124_BO5),
.O6(CLBLM_R_X103Y124_SLICE_X163Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a8080aa0aa000)
  ) CLBLM_R_X103Y124_SLICE_X163Y124_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y124_SLICE_X160Y124_AQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X103Y124_SLICE_X163Y124_DO6),
.I4(CLBLM_L_X98Y122_SLICE_X154Y122_DO6),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y124_SLICE_X163Y124_AO5),
.O6(CLBLM_R_X103Y124_SLICE_X163Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X162Y125_AO5),
.Q(CLBLM_R_X103Y125_SLICE_X162Y125_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X162Y125_CO5),
.Q(CLBLM_R_X103Y125_SLICE_X162Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X162Y125_AO6),
.Q(CLBLM_R_X103Y125_SLICE_X162Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X162Y125_BO6),
.Q(CLBLM_R_X103Y125_SLICE_X162Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X162Y125_CO6),
.Q(CLBLM_R_X103Y125_SLICE_X162Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699696699669)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_DLUT (
.I0(CLBLM_R_X103Y125_SLICE_X162Y125_C5Q),
.I1(CLBLM_R_X103Y125_SLICE_X162Y125_CQ),
.I2(CLBLM_R_X103Y125_SLICE_X163Y125_B5Q),
.I3(CLBLM_R_X103Y125_SLICE_X162Y125_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_DO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y125_SLICE_X162Y125_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X103Y125_SLICE_X162Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_CO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4455445505550555)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_BLUT (
.I0(CLBLM_R_X103Y126_SLICE_X163Y126_CO6),
.I1(CLBLM_R_X103Y125_SLICE_X162Y125_A5Q),
.I2(CLBLM_R_X103Y125_SLICE_X162Y125_DO6),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_BO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X103Y125_SLICE_X162Y125_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y125_SLICE_X162Y125_A5Q),
.I2(CLBLM_R_X103Y123_SLICE_X162Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X162Y125_AO5),
.O6(CLBLM_R_X103Y125_SLICE_X162Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X163Y125_BO5),
.Q(CLBLM_R_X103Y125_SLICE_X163Y125_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X163Y125_CO5),
.Q(CLBLM_R_X103Y125_SLICE_X163Y125_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X163Y125_AO6),
.Q(CLBLM_R_X103Y125_SLICE_X163Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X163Y125_BO6),
.Q(CLBLM_R_X103Y125_SLICE_X163Y125_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y125_SLICE_X163Y125_CO6),
.Q(CLBLM_R_X103Y125_SLICE_X163Y125_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_DLUT (
.I0(CLBLM_R_X103Y125_SLICE_X163Y125_C5Q),
.I1(CLBLM_R_X103Y125_SLICE_X163Y125_CQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y125_SLICE_X163Y125_BQ),
.I4(CLBLM_R_X103Y125_SLICE_X163Y125_AQ),
.I5(RIOB33_X105Y147_IOB_X1Y148_I),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_DO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000c0c0c0c0)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y125_SLICE_X163Y125_CQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X103Y125_SLICE_X163Y125_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_CO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y125_SLICE_X163Y125_AQ),
.I3(CLBLM_R_X103Y125_SLICE_X162Y125_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_BO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ddff11ff)
  ) CLBLM_R_X103Y125_SLICE_X163Y125_ALUT (
.I0(CLBLM_R_X103Y125_SLICE_X163Y125_DO6),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(1'b1),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_R_X103Y125_SLICE_X162Y125_AQ),
.I5(CLBLM_R_X103Y126_SLICE_X163Y126_BO6),
.O5(CLBLM_R_X103Y125_SLICE_X163Y125_AO5),
.O6(CLBLM_R_X103Y125_SLICE_X163Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y126_SLICE_X162Y126_BO5),
.Q(CLBLM_R_X103Y126_SLICE_X162Y126_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y126_SLICE_X162Y126_AO6),
.Q(CLBLM_R_X103Y126_SLICE_X162Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y126_SLICE_X162Y126_BO6),
.Q(CLBLM_R_X103Y126_SLICE_X162Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f066999966)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_DLUT (
.I0(CLBLL_L_X102Y126_SLICE_X161Y126_BQ),
.I1(CLBLM_R_X103Y126_SLICE_X162Y126_AQ),
.I2(CLBLM_R_X101Y126_SLICE_X159Y126_AQ),
.I3(CLBLM_R_X103Y126_SLICE_X162Y126_BQ),
.I4(CLBLM_R_X103Y126_SLICE_X162Y126_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y126_SLICE_X162Y126_DO5),
.O6(CLBLM_R_X103Y126_SLICE_X162Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0069699696)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_CLUT (
.I0(CLBLL_L_X102Y126_SLICE_X161Y126_BQ),
.I1(CLBLM_R_X103Y126_SLICE_X162Y126_AQ),
.I2(CLBLM_R_X103Y126_SLICE_X162Y126_BQ),
.I3(CLBLL_L_X102Y126_SLICE_X161Y126_A5Q),
.I4(CLBLM_R_X103Y126_SLICE_X162Y126_B5Q),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X103Y126_SLICE_X162Y126_CO5),
.O6(CLBLM_R_X103Y126_SLICE_X162Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y126_SLICE_X162Y126_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X102Y126_SLICE_X161Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y126_SLICE_X162Y126_BO5),
.O6(CLBLM_R_X103Y126_SLICE_X162Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa8aaa80008a0080)
  ) CLBLM_R_X103Y126_SLICE_X162Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLL_L_X102Y126_SLICE_X161Y126_DQ),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y119_IOB_X1Y120_I),
.I5(CLBLM_R_X103Y126_SLICE_X162Y126_CO6),
.O5(CLBLM_R_X103Y126_SLICE_X162Y126_AO5),
.O6(CLBLM_R_X103Y126_SLICE_X162Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y126_SLICE_X163Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y126_SLICE_X163Y126_AO5),
.Q(CLBLM_R_X103Y126_SLICE_X163Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y126_SLICE_X163Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y126_SLICE_X163Y126_AO6),
.Q(CLBLM_R_X103Y126_SLICE_X163Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f2f1f3f0f2f1f3f)
  ) CLBLM_R_X103Y126_SLICE_X163Y126_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_B5Q),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y126_SLICE_X163Y126_DO5),
.O6(CLBLM_R_X103Y126_SLICE_X163Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f2f0f2f0f7f0f7f)
  ) CLBLM_R_X103Y126_SLICE_X163Y126_CLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(CLBLM_R_X103Y126_SLICE_X163Y126_AQ),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(1'b1),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X103Y126_SLICE_X163Y126_CO5),
.O6(CLBLM_R_X103Y126_SLICE_X163Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555f55ff555f)
  ) CLBLM_R_X103Y126_SLICE_X163Y126_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(1'b1),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X103Y126_SLICE_X163Y126_A5Q),
.O5(CLBLM_R_X103Y126_SLICE_X163Y126_BO5),
.O6(CLBLM_R_X103Y126_SLICE_X163Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h82828282aa0000aa)
  ) CLBLM_R_X103Y126_SLICE_X163Y126_ALUT (
.I0(RIOB33_X105Y145_IOB_X1Y146_I),
.I1(CLBLM_R_X103Y125_SLICE_X163Y125_B5Q),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_B5Q),
.I3(CLBLM_R_X103Y126_SLICE_X163Y126_AQ),
.I4(CLBLM_R_X103Y125_SLICE_X163Y125_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y126_SLICE_X163Y126_AO5),
.O6(CLBLM_R_X103Y126_SLICE_X163Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y127_SLICE_X162Y127_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.D(CLBLM_R_X103Y127_SLICE_X162Y127_AO6),
.Q(CLBLM_R_X103Y127_SLICE_X162Y127_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X162Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X162Y127_DO5),
.O6(CLBLM_R_X103Y127_SLICE_X162Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X162Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X162Y127_CO5),
.O6(CLBLM_R_X103Y127_SLICE_X162Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X162Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X162Y127_BO5),
.O6(CLBLM_R_X103Y127_SLICE_X162Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccafcca000000000)
  ) CLBLM_R_X103Y127_SLICE_X162Y127_ALUT (
.I0(CLBLL_L_X102Y127_SLICE_X161Y127_B5Q),
.I1(CLBLL_L_X102Y127_SLICE_X161Y127_CO6),
.I2(RIOB33_X105Y147_IOB_X1Y147_I),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(RIOB33_X105Y145_IOB_X1Y146_I),
.O5(CLBLM_R_X103Y127_SLICE_X162Y127_AO5),
.O6(CLBLM_R_X103Y127_SLICE_X162Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X163Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X163Y127_DO5),
.O6(CLBLM_R_X103Y127_SLICE_X163Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X163Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X163Y127_CO5),
.O6(CLBLM_R_X103Y127_SLICE_X163Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X163Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X163Y127_BO5),
.O6(CLBLM_R_X103Y127_SLICE_X163Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y127_SLICE_X163Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y127_SLICE_X163Y127_AO5),
.O6(CLBLM_R_X103Y127_SLICE_X163Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y77_IOB_X1Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y1_IOB_X0Y1_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y1_IOB_X0Y2_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y3_IOB_X0Y3_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y4_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y3_IOB_X0Y4_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y5_IOB_X0Y5_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y5_IOB_X0Y5_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y5_IOB_X0Y6_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y5_IOB_X0Y6_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y51_IOB_X0Y51_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y51_IOB_X0Y51_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y51_IOB_X0Y52_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y51_IOB_X0Y52_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y53_IOB_X0Y53_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y53_IOB_X0Y53_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y53_IOB_X0Y54_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y53_IOB_X0Y54_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y55_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y55_IOB_X0Y55_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y56_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y55_IOB_X0Y56_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y57_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y57_IOB_X0Y57_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y58_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y57_IOB_X0Y58_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y59_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y59_IOB_X0Y59_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y60_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y59_IOB_X0Y60_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y61_IOB_X0Y61_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y61_IOB_X0Y61_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y61_IOB_X0Y62_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y61_IOB_X0Y62_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y63_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y63_IOB_X0Y63_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y67_IOB_X0Y67_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y67_IOB_X0Y67_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y67_IOB_X0Y68_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y67_IOB_X0Y68_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y69_IOB_X0Y69_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y69_IOB_X0Y69_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y69_IOB_X0Y70_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y69_IOB_X0Y70_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y71_IOB_X0Y71_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y71_IOB_X0Y71_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y71_IOB_X0Y72_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y71_IOB_X0Y72_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y73_IOB_X0Y73_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y73_IOB_X0Y73_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y73_IOB_X0Y74_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y73_IOB_X0Y74_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y75_IOB_X0Y75_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y75_IOB_X0Y75_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y75_IOB_X0Y76_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y75_IOB_X0Y76_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y77_IOB_X0Y77_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y77_IOB_X0Y77_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y77_IOB_X0Y78_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y77_IOB_X0Y78_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y79_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y79_IOB_X0Y79_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y81_IOB_X0Y81_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y81_IOB_X0Y81_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y81_IOB_X0Y82_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y81_IOB_X0Y82_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y83_IOB_X0Y83_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y83_IOB_X0Y83_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y83_IOB_X0Y84_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y83_IOB_X0Y84_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y85_IOB_X0Y85_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y85_IOB_X0Y85_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y85_IOB_X0Y86_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y85_IOB_X0Y86_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y87_IOB_X0Y87_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y87_IOB_X0Y87_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y87_IOB_X0Y88_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y87_IOB_X0Y88_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y89_IOB_X0Y89_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y89_IOB_X0Y89_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y89_IOB_X0Y90_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y89_IOB_X0Y90_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y91_IOB_X0Y91_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y91_IOB_X0Y91_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y91_IOB_X0Y92_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y91_IOB_X0Y92_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y93_IOB_X0Y93_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y93_IOB_X0Y93_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y93_IOB_X0Y94_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y93_IOB_X0Y94_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y95_IOB_X0Y95_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y95_IOB_X0Y95_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y95_IOB_X0Y96_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y95_IOB_X0Y96_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y97_IOB_X0Y97_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y97_IOB_X0Y97_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y97_IOB_X0Y98_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y97_IOB_X0Y98_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y201_IOB_X0Y201_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y201_IOB_X0Y201_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y201_IOB_X0Y202_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y201_IOB_X0Y202_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y203_IOB_X0Y203_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y203_IOB_X0Y203_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y203_IOB_X0Y204_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y203_IOB_X0Y204_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y205_IOB_X0Y205_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y205_IOB_X0Y205_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y205_IOB_X0Y206_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y205_IOB_X0Y206_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y207_IOB_X0Y207_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y207_IOB_X0Y207_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y207_IOB_X0Y208_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y207_IOB_X0Y208_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y209_IOB_X0Y209_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y209_IOB_X0Y209_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y209_IOB_X0Y210_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y209_IOB_X0Y210_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y211_IOB_X0Y211_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y211_IOB_X0Y211_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y211_IOB_X0Y212_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y211_IOB_X0Y212_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y213_IOB_X0Y213_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y213_IOB_X0Y213_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y213_IOB_X0Y214_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y213_IOB_X0Y214_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y215_IOB_X0Y215_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y215_IOB_X0Y215_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y215_IOB_X0Y216_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y215_IOB_X0Y216_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y217_IOB_X0Y217_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y217_IOB_X0Y217_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y217_IOB_X0Y218_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y217_IOB_X0Y218_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y219_IOB_X0Y219_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y219_IOB_X0Y219_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y219_IOB_X0Y220_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y219_IOB_X0Y220_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y221_IOB_X0Y221_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y221_IOB_X0Y221_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y221_IOB_X0Y222_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y221_IOB_X0Y222_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y223_IOB_X0Y223_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y223_IOB_X0Y223_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y223_IOB_X0Y224_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y223_IOB_X0Y224_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y225_IOB_X0Y225_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y225_IOB_X0Y225_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y225_IOB_X0Y226_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y225_IOB_X0Y226_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y227_IOB_X0Y227_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y227_IOB_X0Y227_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y227_IOB_X0Y228_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y227_IOB_X0Y228_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y229_IOB_X0Y229_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y229_IOB_X0Y229_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y229_IOB_X0Y230_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y229_IOB_X0Y230_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y231_IOB_X0Y231_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y231_IOB_X0Y231_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y231_IOB_X0Y232_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y231_IOB_X0Y232_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y233_IOB_X0Y233_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y233_IOB_X0Y233_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y233_IOB_X0Y234_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y233_IOB_X0Y234_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y235_IOB_X0Y235_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y235_IOB_X0Y235_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y235_IOB_X0Y236_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y235_IOB_X0Y236_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y237_IOB_X0Y237_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y237_IOB_X0Y237_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y237_IOB_X0Y238_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y237_IOB_X0Y238_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y239_IOB_X0Y239_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y239_IOB_X0Y239_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y239_IOB_X0Y240_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y239_IOB_X0Y240_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y241_IOB_X0Y241_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y241_IOB_X0Y241_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y241_IOB_X0Y242_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y241_IOB_X0Y242_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y243_IOB_X0Y243_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y243_IOB_X0Y243_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y243_IOB_X0Y244_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y243_IOB_X0Y244_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y245_IOB_X0Y245_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y245_IOB_X0Y245_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y245_IOB_X0Y246_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y245_IOB_X0Y246_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y247_IOB_X0Y247_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y247_IOB_X0Y247_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_X0Y247_IOB_X0Y248_OBUFT (
.I(1'b0),
.O(LIOB33_X0Y247_IOB_X0Y248_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y0_IOB_X0Y0_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y50_IOB_X0Y50_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y99_IOB_X0Y99_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y200_IOB_X0Y200_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y200_IOB_X0Y200_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y249_IOB_X0Y249_OBUFT (
.I(1'b0),
.O(LIOB33_SING_X0Y249_IOB_X0Y249_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y51_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y51_IOB_X1Y51_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y52_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y51_IOB_X1Y52_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y53_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y53_IOB_X1Y53_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y54_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y53_IOB_X1Y54_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y55_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y55_IOB_X1Y55_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y56_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y55_IOB_X1Y56_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y57_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y57_IOB_X1Y57_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y58_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y57_IOB_X1Y58_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y59_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y59_IOB_X1Y59_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y60_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y59_IOB_X1Y60_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y61_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y61_IOB_X1Y61_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y62_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y61_IOB_X1Y62_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y63_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y63_IOB_X1Y63_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y64_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y63_IOB_X1Y64_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y65_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y65_IOB_X1Y65_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y66_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y65_IOB_X1Y66_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y67_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y67_IOB_X1Y67_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y68_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y67_IOB_X1Y68_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y69_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y69_IOB_X1Y69_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y70_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y69_IOB_X1Y70_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y71_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y71_IOB_X1Y71_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y72_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y71_IOB_X1Y72_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y73_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y73_IOB_X1Y73_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y74_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y73_IOB_X1Y74_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y75_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y75_IOB_X1Y75_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y76_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y75_IOB_X1Y76_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y77_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y77_IOB_X1Y77_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y77_IOB_X1Y78_IBUF (
.I(RIOB33_X105Y77_IOB_X1Y78_IPAD),
.O(RIOB33_X105Y77_IOB_X1Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y79_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y79_IOB_X1Y79_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y80_OBUF (
.I(CLBLM_R_X103Y119_SLICE_X163Y119_CO6),
.O(RIOB33_X105Y79_IOB_X1Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y81_OBUF (
.I(CLBLL_L_X102Y119_SLICE_X161Y119_CO6),
.O(RIOB33_X105Y81_IOB_X1Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y82_OBUF (
.I(CLBLM_R_X101Y120_SLICE_X159Y120_CO6),
.O(RIOB33_X105Y81_IOB_X1Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y83_OBUF (
.I(CLBLL_L_X102Y117_SLICE_X160Y117_CO6),
.O(RIOB33_X105Y83_IOB_X1Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y84_OBUF (
.I(CLBLM_R_X101Y119_SLICE_X159Y119_CO6),
.O(RIOB33_X105Y83_IOB_X1Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y85_OBUF (
.I(CLBLM_R_X103Y116_SLICE_X162Y116_CO6),
.O(RIOB33_X105Y85_IOB_X1Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y86_OBUF (
.I(CLBLM_R_X103Y117_SLICE_X162Y117_CO6),
.O(RIOB33_X105Y85_IOB_X1Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y87_OBUF (
.I(CLBLL_L_X100Y115_SLICE_X157Y115_CO6),
.O(RIOB33_X105Y87_IOB_X1Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y88_OBUF (
.I(CLBLM_R_X101Y117_SLICE_X159Y117_AO5),
.O(RIOB33_X105Y87_IOB_X1Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y89_OBUF (
.I(CLBLM_R_X101Y116_SLICE_X159Y116_AO6),
.O(RIOB33_X105Y89_IOB_X1Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y90_OBUF (
.I(CLBLL_L_X102Y116_SLICE_X160Y116_AO6),
.O(RIOB33_X105Y89_IOB_X1Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y91_OBUF (
.I(CLBLL_L_X102Y115_SLICE_X161Y115_AO6),
.O(RIOB33_X105Y91_IOB_X1Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y92_OBUF (
.I(CLBLL_L_X102Y119_SLICE_X160Y119_CO6),
.O(RIOB33_X105Y91_IOB_X1Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y93_OBUF (
.I(CLBLL_L_X102Y114_SLICE_X160Y114_AO6),
.O(RIOB33_X105Y93_IOB_X1Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y94_OBUF (
.I(CLBLM_R_X103Y113_SLICE_X163Y113_AO6),
.O(RIOB33_X105Y93_IOB_X1Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y95_OBUF (
.I(CLBLM_R_X103Y113_SLICE_X163Y113_BO6),
.O(RIOB33_X105Y95_IOB_X1Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y96_OBUF (
.I(CLBLM_R_X103Y112_SLICE_X162Y112_AO6),
.O(RIOB33_X105Y95_IOB_X1Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y97_OBUF (
.I(CLBLM_R_X103Y111_SLICE_X162Y111_AO6),
.O(RIOB33_X105Y97_IOB_X1Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y98_OBUF (
.I(CLBLL_L_X102Y111_SLICE_X161Y111_AO6),
.O(RIOB33_X105Y97_IOB_X1Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y101_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y101_IOB_X1Y101_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y102_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y101_IOB_X1Y102_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y103_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y103_IOB_X1Y103_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y104_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y103_IOB_X1Y104_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y105_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y105_IOB_X1Y105_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y106_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y105_IOB_X1Y106_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(CLBLL_L_X102Y112_SLICE_X160Y112_AO6),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(CLBLM_R_X101Y113_SLICE_X159Y113_AO6),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(CLBLM_R_X101Y113_SLICE_X159Y113_BO6),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLM_R_X103Y121_SLICE_X162Y121_CO6),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLM_R_X101Y116_SLICE_X159Y116_BO6),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUFT (
.I(1'b0),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLL_L_X102Y118_SLICE_X160Y118_AO6),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X103Y120_SLICE_X163Y120_CO6),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLL_L_X102Y120_SLICE_X161Y120_CO6),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_R_X103Y124_SLICE_X162Y124_CO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLL_L_X102Y124_SLICE_X161Y124_CO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X103Y124_SLICE_X163Y124_CO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y50_IOB_X1Y50_OBUFT (
.I(1'b0),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y99_IOB_X1Y99_OBUF (
.I(CLBLL_L_X102Y111_SLICE_X160Y111_AO6),
.O(RIOB33_SING_X105Y99_IOB_X1Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_OBUFT (
.I(1'b0),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUFT #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUFT (
.I(1'b0),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD),
.T(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLL_L_X102Y123_SLICE_X160Y123_CO6),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A = CLBLL_L_X100Y111_SLICE_X156Y111_AO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B = CLBLL_L_X100Y111_SLICE_X156Y111_BO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C = CLBLL_L_X100Y111_SLICE_X156Y111_CO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D = CLBLL_L_X100Y111_SLICE_X156Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_AMUX = CLBLL_L_X100Y111_SLICE_X156Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_BMUX = CLBLL_L_X100Y111_SLICE_X156Y111_B5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A = CLBLL_L_X100Y111_SLICE_X157Y111_AO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B = CLBLL_L_X100Y111_SLICE_X157Y111_BO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C = CLBLL_L_X100Y111_SLICE_X157Y111_CO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D = CLBLL_L_X100Y111_SLICE_X157Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_AMUX = CLBLL_L_X100Y111_SLICE_X157Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_BMUX = CLBLL_L_X100Y111_SLICE_X157Y111_B5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_CMUX = CLBLL_L_X100Y111_SLICE_X157Y111_C5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_DMUX = CLBLL_L_X100Y111_SLICE_X157Y111_DO6;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A = CLBLL_L_X100Y112_SLICE_X156Y112_AO6;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B = CLBLL_L_X100Y112_SLICE_X156Y112_BO6;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C = CLBLL_L_X100Y112_SLICE_X156Y112_CO6;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D = CLBLL_L_X100Y112_SLICE_X156Y112_DO6;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_AMUX = CLBLL_L_X100Y112_SLICE_X156Y112_A5Q;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A = CLBLL_L_X100Y112_SLICE_X157Y112_AO6;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B = CLBLL_L_X100Y112_SLICE_X157Y112_BO6;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C = CLBLL_L_X100Y112_SLICE_X157Y112_CO6;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D = CLBLL_L_X100Y112_SLICE_X157Y112_DO6;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_AMUX = CLBLL_L_X100Y112_SLICE_X157Y112_A5Q;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A = CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B = CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C = CLBLL_L_X100Y113_SLICE_X156Y113_CO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D = CLBLL_L_X100Y113_SLICE_X156Y113_DO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_AMUX = CLBLL_L_X100Y113_SLICE_X156Y113_A5Q;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_BMUX = CLBLL_L_X100Y113_SLICE_X156Y113_B5Q;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_CMUX = CLBLL_L_X100Y113_SLICE_X156Y113_C5Q;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A = CLBLL_L_X100Y113_SLICE_X157Y113_AO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B = CLBLL_L_X100Y113_SLICE_X157Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C = CLBLL_L_X100Y113_SLICE_X157Y113_CO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D = CLBLL_L_X100Y113_SLICE_X157Y113_DO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_AMUX = CLBLL_L_X100Y113_SLICE_X157Y113_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A = CLBLL_L_X100Y114_SLICE_X156Y114_AO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B = CLBLL_L_X100Y114_SLICE_X156Y114_BO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C = CLBLL_L_X100Y114_SLICE_X156Y114_CO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D = CLBLL_L_X100Y114_SLICE_X156Y114_DO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_AMUX = CLBLL_L_X100Y114_SLICE_X156Y114_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_BMUX = CLBLL_L_X100Y114_SLICE_X156Y114_B5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_DMUX = CLBLL_L_X100Y114_SLICE_X156Y114_DO6;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A = CLBLL_L_X100Y114_SLICE_X157Y114_AO6;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B = CLBLL_L_X100Y114_SLICE_X157Y114_BO6;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C = CLBLL_L_X100Y114_SLICE_X157Y114_CO6;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D = CLBLL_L_X100Y114_SLICE_X157Y114_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A = CLBLL_L_X100Y115_SLICE_X156Y115_AO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B = CLBLL_L_X100Y115_SLICE_X156Y115_BO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C = CLBLL_L_X100Y115_SLICE_X156Y115_CO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D = CLBLL_L_X100Y115_SLICE_X156Y115_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_AMUX = CLBLL_L_X100Y115_SLICE_X156Y115_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_BMUX = CLBLL_L_X100Y115_SLICE_X156Y115_B5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_CMUX = CLBLL_L_X100Y115_SLICE_X156Y115_C5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A = CLBLL_L_X100Y115_SLICE_X157Y115_AO6;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B = CLBLL_L_X100Y115_SLICE_X157Y115_BO6;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C = CLBLL_L_X100Y115_SLICE_X157Y115_CO6;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D = CLBLL_L_X100Y115_SLICE_X157Y115_DO6;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_BMUX = CLBLL_L_X100Y115_SLICE_X157Y115_B5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_DMUX = CLBLL_L_X100Y115_SLICE_X157Y115_DO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A = CLBLL_L_X100Y116_SLICE_X156Y116_AO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B = CLBLL_L_X100Y116_SLICE_X156Y116_BO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C = CLBLL_L_X100Y116_SLICE_X156Y116_CO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D = CLBLL_L_X100Y116_SLICE_X156Y116_DO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_AMUX = CLBLL_L_X100Y116_SLICE_X156Y116_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_BMUX = CLBLL_L_X100Y116_SLICE_X156Y116_B5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_CMUX = CLBLL_L_X100Y116_SLICE_X156Y116_CO6;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A = CLBLL_L_X100Y116_SLICE_X157Y116_AO6;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B = CLBLL_L_X100Y116_SLICE_X157Y116_BO6;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C = CLBLL_L_X100Y116_SLICE_X157Y116_CO6;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D = CLBLL_L_X100Y116_SLICE_X157Y116_DO6;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_AMUX = CLBLL_L_X100Y116_SLICE_X157Y116_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_BMUX = CLBLL_L_X100Y116_SLICE_X157Y116_B5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A = CLBLL_L_X100Y117_SLICE_X156Y117_AO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B = CLBLL_L_X100Y117_SLICE_X156Y117_BO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C = CLBLL_L_X100Y117_SLICE_X156Y117_CO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D = CLBLL_L_X100Y117_SLICE_X156Y117_DO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_AMUX = CLBLL_L_X100Y117_SLICE_X156Y117_A5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_BMUX = CLBLL_L_X100Y117_SLICE_X156Y117_B5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_CMUX = CLBLL_L_X100Y117_SLICE_X156Y117_CO6;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A = CLBLL_L_X100Y117_SLICE_X157Y117_AO6;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B = CLBLL_L_X100Y117_SLICE_X157Y117_BO6;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C = CLBLL_L_X100Y117_SLICE_X157Y117_CO6;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D = CLBLL_L_X100Y117_SLICE_X157Y117_DO6;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_AMUX = CLBLL_L_X100Y117_SLICE_X157Y117_A5Q;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_BMUX = CLBLL_L_X100Y117_SLICE_X157Y117_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A = CLBLL_L_X100Y118_SLICE_X156Y118_AO6;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B = CLBLL_L_X100Y118_SLICE_X156Y118_BO6;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C = CLBLL_L_X100Y118_SLICE_X156Y118_CO6;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D = CLBLL_L_X100Y118_SLICE_X156Y118_DO6;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_AMUX = CLBLL_L_X100Y118_SLICE_X156Y118_A5Q;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_BMUX = CLBLL_L_X100Y118_SLICE_X156Y118_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A = CLBLL_L_X100Y118_SLICE_X157Y118_AO6;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B = CLBLL_L_X100Y118_SLICE_X157Y118_BO6;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C = CLBLL_L_X100Y118_SLICE_X157Y118_CO6;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D = CLBLL_L_X100Y118_SLICE_X157Y118_DO6;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_AMUX = CLBLL_L_X100Y118_SLICE_X157Y118_A5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_BMUX = CLBLL_L_X100Y118_SLICE_X157Y118_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_CMUX = CLBLL_L_X100Y118_SLICE_X157Y118_C5Q;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A = CLBLL_L_X100Y119_SLICE_X156Y119_AO6;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B = CLBLL_L_X100Y119_SLICE_X156Y119_BO6;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C = CLBLL_L_X100Y119_SLICE_X156Y119_CO6;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D = CLBLL_L_X100Y119_SLICE_X156Y119_DO6;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_BMUX = CLBLL_L_X100Y119_SLICE_X156Y119_B5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A = CLBLL_L_X100Y119_SLICE_X157Y119_AO6;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B = CLBLL_L_X100Y119_SLICE_X157Y119_BO6;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C = CLBLL_L_X100Y119_SLICE_X157Y119_CO6;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D = CLBLL_L_X100Y119_SLICE_X157Y119_DO6;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_AMUX = CLBLL_L_X100Y119_SLICE_X157Y119_A5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_BMUX = CLBLL_L_X100Y119_SLICE_X157Y119_BO5;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_CMUX = CLBLL_L_X100Y119_SLICE_X157Y119_C5Q;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A = CLBLL_L_X100Y120_SLICE_X156Y120_AO6;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B = CLBLL_L_X100Y120_SLICE_X156Y120_BO6;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C = CLBLL_L_X100Y120_SLICE_X156Y120_CO6;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D = CLBLL_L_X100Y120_SLICE_X156Y120_DO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A = CLBLL_L_X100Y120_SLICE_X157Y120_AO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B = CLBLL_L_X100Y120_SLICE_X157Y120_BO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C = CLBLL_L_X100Y120_SLICE_X157Y120_CO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D = CLBLL_L_X100Y120_SLICE_X157Y120_DO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_AMUX = CLBLL_L_X100Y120_SLICE_X157Y120_A5Q;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A = CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B = CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C = CLBLL_L_X100Y121_SLICE_X156Y121_CO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D = CLBLL_L_X100Y121_SLICE_X156Y121_DO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_AMUX = CLBLL_L_X100Y121_SLICE_X156Y121_A5Q;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_CMUX = CLBLL_L_X100Y121_SLICE_X156Y121_C5Q;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A = CLBLL_L_X100Y121_SLICE_X157Y121_AO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B = CLBLL_L_X100Y121_SLICE_X157Y121_BO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C = CLBLL_L_X100Y121_SLICE_X157Y121_CO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D = CLBLL_L_X100Y121_SLICE_X157Y121_DO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_CMUX = CLBLL_L_X100Y121_SLICE_X157Y121_C5Q;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A = CLBLL_L_X100Y122_SLICE_X156Y122_AO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B = CLBLL_L_X100Y122_SLICE_X156Y122_BO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C = CLBLL_L_X100Y122_SLICE_X156Y122_CO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D = CLBLL_L_X100Y122_SLICE_X156Y122_DO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_AMUX = CLBLL_L_X100Y122_SLICE_X156Y122_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A = CLBLL_L_X100Y122_SLICE_X157Y122_AO6;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B = CLBLL_L_X100Y122_SLICE_X157Y122_BO6;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C = CLBLL_L_X100Y122_SLICE_X157Y122_CO6;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D = CLBLL_L_X100Y122_SLICE_X157Y122_DO6;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_AMUX = CLBLL_L_X100Y122_SLICE_X157Y122_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_BMUX = CLBLL_L_X100Y122_SLICE_X157Y122_B5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_CMUX = CLBLL_L_X100Y122_SLICE_X157Y122_C5Q;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A = CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B = CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C = CLBLL_L_X100Y123_SLICE_X156Y123_CO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D = CLBLL_L_X100Y123_SLICE_X156Y123_DO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_AMUX = CLBLL_L_X100Y123_SLICE_X156Y123_A5Q;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_BMUX = CLBLL_L_X100Y123_SLICE_X156Y123_B5Q;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A = CLBLL_L_X100Y123_SLICE_X157Y123_AO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B = CLBLL_L_X100Y123_SLICE_X157Y123_BO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C = CLBLL_L_X100Y123_SLICE_X157Y123_CO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D = CLBLL_L_X100Y123_SLICE_X157Y123_DO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_AMUX = CLBLL_L_X100Y123_SLICE_X157Y123_A5Q;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A = CLBLL_L_X100Y124_SLICE_X156Y124_AO6;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B = CLBLL_L_X100Y124_SLICE_X156Y124_BO6;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C = CLBLL_L_X100Y124_SLICE_X156Y124_CO6;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D = CLBLL_L_X100Y124_SLICE_X156Y124_DO6;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_AMUX = CLBLL_L_X100Y124_SLICE_X156Y124_AO6;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_BMUX = CLBLL_L_X100Y124_SLICE_X156Y124_B5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A = CLBLL_L_X100Y124_SLICE_X157Y124_AO6;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B = CLBLL_L_X100Y124_SLICE_X157Y124_BO6;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C = CLBLL_L_X100Y124_SLICE_X157Y124_CO6;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D = CLBLL_L_X100Y124_SLICE_X157Y124_DO6;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_AMUX = CLBLL_L_X100Y124_SLICE_X157Y124_A5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_BMUX = CLBLL_L_X100Y124_SLICE_X157Y124_B5Q;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A = CLBLL_L_X100Y125_SLICE_X156Y125_AO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B = CLBLL_L_X100Y125_SLICE_X156Y125_BO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C = CLBLL_L_X100Y125_SLICE_X156Y125_CO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D = CLBLL_L_X100Y125_SLICE_X156Y125_DO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_BMUX = CLBLL_L_X100Y125_SLICE_X156Y125_B5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A = CLBLL_L_X100Y125_SLICE_X157Y125_AO6;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B = CLBLL_L_X100Y125_SLICE_X157Y125_BO6;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C = CLBLL_L_X100Y125_SLICE_X157Y125_CO6;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D = CLBLL_L_X100Y125_SLICE_X157Y125_DO6;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_AMUX = CLBLL_L_X100Y125_SLICE_X157Y125_A5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_BMUX = CLBLL_L_X100Y125_SLICE_X157Y125_B5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_CMUX = CLBLL_L_X100Y125_SLICE_X157Y125_C5Q;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A = CLBLL_L_X100Y126_SLICE_X156Y126_AO6;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B = CLBLL_L_X100Y126_SLICE_X156Y126_BO6;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C = CLBLL_L_X100Y126_SLICE_X156Y126_CO6;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D = CLBLL_L_X100Y126_SLICE_X156Y126_DO6;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_AMUX = CLBLL_L_X100Y126_SLICE_X156Y126_A5Q;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_BMUX = CLBLL_L_X100Y126_SLICE_X156Y126_B5Q;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_CMUX = CLBLL_L_X100Y126_SLICE_X156Y126_CO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A = CLBLL_L_X100Y126_SLICE_X157Y126_AO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B = CLBLL_L_X100Y126_SLICE_X157Y126_BO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C = CLBLL_L_X100Y126_SLICE_X157Y126_CO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D = CLBLL_L_X100Y126_SLICE_X157Y126_DO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_AMUX = CLBLL_L_X100Y126_SLICE_X157Y126_A5Q;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A = CLBLL_L_X100Y127_SLICE_X156Y127_AO6;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B = CLBLL_L_X100Y127_SLICE_X156Y127_BO6;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C = CLBLL_L_X100Y127_SLICE_X156Y127_CO6;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D = CLBLL_L_X100Y127_SLICE_X156Y127_DO6;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_AMUX = CLBLL_L_X100Y127_SLICE_X156Y127_A5Q;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_BMUX = CLBLL_L_X100Y127_SLICE_X156Y127_B5Q;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A = CLBLL_L_X100Y127_SLICE_X157Y127_AO6;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B = CLBLL_L_X100Y127_SLICE_X157Y127_BO6;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C = CLBLL_L_X100Y127_SLICE_X157Y127_CO6;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D = CLBLL_L_X100Y127_SLICE_X157Y127_DO6;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_BMUX = CLBLL_L_X100Y127_SLICE_X157Y127_B5Q;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A = CLBLL_L_X100Y128_SLICE_X156Y128_AO6;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B = CLBLL_L_X100Y128_SLICE_X156Y128_BO6;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C = CLBLL_L_X100Y128_SLICE_X156Y128_CO6;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D = CLBLL_L_X100Y128_SLICE_X156Y128_DO6;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_AMUX = CLBLL_L_X100Y128_SLICE_X156Y128_A5Q;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A = CLBLL_L_X100Y128_SLICE_X157Y128_AO6;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B = CLBLL_L_X100Y128_SLICE_X157Y128_BO6;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C = CLBLL_L_X100Y128_SLICE_X157Y128_CO6;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D = CLBLL_L_X100Y128_SLICE_X157Y128_DO6;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A = CLBLL_L_X100Y129_SLICE_X156Y129_AO6;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B = CLBLL_L_X100Y129_SLICE_X156Y129_BO6;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C = CLBLL_L_X100Y129_SLICE_X156Y129_CO6;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D = CLBLL_L_X100Y129_SLICE_X156Y129_DO6;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A = CLBLL_L_X100Y129_SLICE_X157Y129_AO6;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B = CLBLL_L_X100Y129_SLICE_X157Y129_BO6;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C = CLBLL_L_X100Y129_SLICE_X157Y129_CO6;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D = CLBLL_L_X100Y129_SLICE_X157Y129_DO6;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_AMUX = CLBLL_L_X100Y129_SLICE_X157Y129_A5Q;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A = CLBLL_L_X100Y130_SLICE_X156Y130_AO6;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B = CLBLL_L_X100Y130_SLICE_X156Y130_BO6;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C = CLBLL_L_X100Y130_SLICE_X156Y130_CO6;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D = CLBLL_L_X100Y130_SLICE_X156Y130_DO6;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A = CLBLL_L_X100Y130_SLICE_X157Y130_AO6;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B = CLBLL_L_X100Y130_SLICE_X157Y130_BO6;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C = CLBLL_L_X100Y130_SLICE_X157Y130_CO6;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D = CLBLL_L_X100Y130_SLICE_X157Y130_DO6;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A = CLBLL_L_X100Y133_SLICE_X156Y133_AO6;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B = CLBLL_L_X100Y133_SLICE_X156Y133_BO6;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C = CLBLL_L_X100Y133_SLICE_X156Y133_CO6;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D = CLBLL_L_X100Y133_SLICE_X156Y133_DO6;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_AMUX = CLBLL_L_X100Y133_SLICE_X156Y133_A5Q;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A = CLBLL_L_X100Y133_SLICE_X157Y133_AO6;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B = CLBLL_L_X100Y133_SLICE_X157Y133_BO6;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C = CLBLL_L_X100Y133_SLICE_X157Y133_CO6;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D = CLBLL_L_X100Y133_SLICE_X157Y133_DO6;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A = CLBLL_L_X100Y134_SLICE_X156Y134_AO6;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B = CLBLL_L_X100Y134_SLICE_X156Y134_BO6;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C = CLBLL_L_X100Y134_SLICE_X156Y134_CO6;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D = CLBLL_L_X100Y134_SLICE_X156Y134_DO6;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_AMUX = CLBLL_L_X100Y134_SLICE_X156Y134_A5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_BMUX = CLBLL_L_X100Y134_SLICE_X156Y134_B5Q;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A = CLBLL_L_X100Y134_SLICE_X157Y134_AO6;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B = CLBLL_L_X100Y134_SLICE_X157Y134_BO6;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C = CLBLL_L_X100Y134_SLICE_X157Y134_CO6;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D = CLBLL_L_X100Y134_SLICE_X157Y134_DO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A = CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B = CLBLL_L_X102Y111_SLICE_X160Y111_BO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C = CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_AMUX = CLBLL_L_X102Y111_SLICE_X160Y111_AO5;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_BMUX = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_CMUX = CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_DMUX = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A = CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B = CLBLL_L_X102Y111_SLICE_X161Y111_BO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C = CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D = CLBLL_L_X102Y111_SLICE_X161Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_BMUX = CLBLL_L_X102Y111_SLICE_X161Y111_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_CMUX = CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A = CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B = CLBLL_L_X102Y112_SLICE_X160Y112_BO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C = CLBLL_L_X102Y112_SLICE_X160Y112_CO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D = CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_BMUX = CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_DMUX = CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A = CLBLL_L_X102Y112_SLICE_X161Y112_AO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B = CLBLL_L_X102Y112_SLICE_X161Y112_BO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D = CLBLL_L_X102Y112_SLICE_X161Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_AMUX = CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_BMUX = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_CMUX = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A = CLBLL_L_X102Y113_SLICE_X160Y113_AO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B = CLBLL_L_X102Y113_SLICE_X160Y113_BO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C = CLBLL_L_X102Y113_SLICE_X160Y113_CO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D = CLBLL_L_X102Y113_SLICE_X160Y113_DO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_AMUX = CLBLL_L_X102Y113_SLICE_X160Y113_A5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A = CLBLL_L_X102Y113_SLICE_X161Y113_AO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B = CLBLL_L_X102Y113_SLICE_X161Y113_BO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C = CLBLL_L_X102Y113_SLICE_X161Y113_CO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D = CLBLL_L_X102Y113_SLICE_X161Y113_DO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_AMUX = CLBLL_L_X102Y113_SLICE_X161Y113_A5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_BMUX = CLBLL_L_X102Y113_SLICE_X161Y113_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_CMUX = CLBLL_L_X102Y113_SLICE_X161Y113_CO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A = CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B = CLBLL_L_X102Y114_SLICE_X160Y114_BO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C = CLBLL_L_X102Y114_SLICE_X160Y114_CO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D = CLBLL_L_X102Y114_SLICE_X160Y114_DO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_AMUX = CLBLL_L_X102Y114_SLICE_X160Y114_AO5;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_BMUX = CLBLL_L_X102Y114_SLICE_X160Y114_B5Q;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_CMUX = CLBLL_L_X102Y114_SLICE_X160Y114_C5Q;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A = CLBLL_L_X102Y114_SLICE_X161Y114_AO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B = CLBLL_L_X102Y114_SLICE_X161Y114_BO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C = CLBLL_L_X102Y114_SLICE_X161Y114_CO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D = CLBLL_L_X102Y114_SLICE_X161Y114_DO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_AMUX = CLBLL_L_X102Y114_SLICE_X161Y114_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A = CLBLL_L_X102Y115_SLICE_X160Y115_AO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B = CLBLL_L_X102Y115_SLICE_X160Y115_BO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C = CLBLL_L_X102Y115_SLICE_X160Y115_CO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D = CLBLL_L_X102Y115_SLICE_X160Y115_DO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_AMUX = CLBLL_L_X102Y115_SLICE_X160Y115_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_BMUX = CLBLL_L_X102Y115_SLICE_X160Y115_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_CMUX = CLBLL_L_X102Y115_SLICE_X160Y115_CO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A = CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B = CLBLL_L_X102Y115_SLICE_X161Y115_BO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C = CLBLL_L_X102Y115_SLICE_X161Y115_CO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D = CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_AMUX = CLBLL_L_X102Y115_SLICE_X161Y115_AO5;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_BMUX = CLBLL_L_X102Y115_SLICE_X161Y115_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_CMUX = CLBLL_L_X102Y115_SLICE_X161Y115_C5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A = CLBLL_L_X102Y116_SLICE_X160Y116_AO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B = CLBLL_L_X102Y116_SLICE_X160Y116_BO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C = CLBLL_L_X102Y116_SLICE_X160Y116_CO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D = CLBLL_L_X102Y116_SLICE_X160Y116_DO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_AMUX = CLBLL_L_X102Y116_SLICE_X160Y116_AO5;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_BMUX = CLBLL_L_X102Y116_SLICE_X160Y116_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_CMUX = CLBLL_L_X102Y116_SLICE_X160Y116_C5Q;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A = CLBLL_L_X102Y116_SLICE_X161Y116_AO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B = CLBLL_L_X102Y116_SLICE_X161Y116_BO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C = CLBLL_L_X102Y116_SLICE_X161Y116_CO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D = CLBLL_L_X102Y116_SLICE_X161Y116_DO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_AMUX = CLBLL_L_X102Y116_SLICE_X161Y116_A5Q;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_BMUX = CLBLL_L_X102Y116_SLICE_X161Y116_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_CMUX = CLBLL_L_X102Y116_SLICE_X161Y116_CO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_DMUX = CLBLL_L_X102Y116_SLICE_X161Y116_DO6;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A = CLBLL_L_X102Y117_SLICE_X160Y117_AO6;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B = CLBLL_L_X102Y117_SLICE_X160Y117_BO6;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C = CLBLL_L_X102Y117_SLICE_X160Y117_CO6;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D = CLBLL_L_X102Y117_SLICE_X160Y117_DO6;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_BMUX = CLBLL_L_X102Y117_SLICE_X160Y117_B5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A = CLBLL_L_X102Y117_SLICE_X161Y117_AO6;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B = CLBLL_L_X102Y117_SLICE_X161Y117_BO6;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C = CLBLL_L_X102Y117_SLICE_X161Y117_CO6;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D = CLBLL_L_X102Y117_SLICE_X161Y117_DO6;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_AMUX = CLBLL_L_X102Y117_SLICE_X161Y117_A5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_BMUX = CLBLL_L_X102Y117_SLICE_X161Y117_B5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_CMUX = CLBLL_L_X102Y117_SLICE_X161Y117_C5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_DMUX = CLBLL_L_X102Y117_SLICE_X161Y117_D5Q;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A = CLBLL_L_X102Y118_SLICE_X160Y118_AO6;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B = CLBLL_L_X102Y118_SLICE_X160Y118_BO6;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C = CLBLL_L_X102Y118_SLICE_X160Y118_CO6;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D = CLBLL_L_X102Y118_SLICE_X160Y118_DO6;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_AMUX = CLBLL_L_X102Y118_SLICE_X160Y118_AO5;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A = CLBLL_L_X102Y118_SLICE_X161Y118_AO6;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B = CLBLL_L_X102Y118_SLICE_X161Y118_BO6;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C = CLBLL_L_X102Y118_SLICE_X161Y118_CO6;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D = CLBLL_L_X102Y118_SLICE_X161Y118_DO6;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A = CLBLL_L_X102Y119_SLICE_X160Y119_AO6;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B = CLBLL_L_X102Y119_SLICE_X160Y119_BO6;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C = CLBLL_L_X102Y119_SLICE_X160Y119_CO6;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D = CLBLL_L_X102Y119_SLICE_X160Y119_DO6;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_AMUX = CLBLL_L_X102Y119_SLICE_X160Y119_A5Q;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_BMUX = CLBLL_L_X102Y119_SLICE_X160Y119_B5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A = CLBLL_L_X102Y119_SLICE_X161Y119_AO6;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B = CLBLL_L_X102Y119_SLICE_X161Y119_BO6;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C = CLBLL_L_X102Y119_SLICE_X161Y119_CO6;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D = CLBLL_L_X102Y119_SLICE_X161Y119_DO6;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_BMUX = CLBLL_L_X102Y119_SLICE_X161Y119_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A = CLBLL_L_X102Y120_SLICE_X160Y120_AO6;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B = CLBLL_L_X102Y120_SLICE_X160Y120_BO6;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C = CLBLL_L_X102Y120_SLICE_X160Y120_CO6;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D = CLBLL_L_X102Y120_SLICE_X160Y120_DO6;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_BMUX = CLBLL_L_X102Y120_SLICE_X160Y120_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_CMUX = CLBLL_L_X102Y120_SLICE_X160Y120_C5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_DMUX = CLBLL_L_X102Y120_SLICE_X160Y120_D5Q;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A = CLBLL_L_X102Y120_SLICE_X161Y120_AO6;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B = CLBLL_L_X102Y120_SLICE_X161Y120_BO6;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C = CLBLL_L_X102Y120_SLICE_X161Y120_CO6;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D = CLBLL_L_X102Y120_SLICE_X161Y120_DO6;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_BMUX = CLBLL_L_X102Y120_SLICE_X161Y120_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_DMUX = CLBLL_L_X102Y120_SLICE_X161Y120_DO6;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A = CLBLL_L_X102Y121_SLICE_X160Y121_AO6;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B = CLBLL_L_X102Y121_SLICE_X160Y121_BO6;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C = CLBLL_L_X102Y121_SLICE_X160Y121_CO6;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D = CLBLL_L_X102Y121_SLICE_X160Y121_DO6;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A = CLBLL_L_X102Y121_SLICE_X161Y121_AO6;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B = CLBLL_L_X102Y121_SLICE_X161Y121_BO6;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C = CLBLL_L_X102Y121_SLICE_X161Y121_CO6;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D = CLBLL_L_X102Y121_SLICE_X161Y121_DO6;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_AMUX = CLBLL_L_X102Y121_SLICE_X161Y121_A5Q;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_BMUX = CLBLL_L_X102Y121_SLICE_X161Y121_B5Q;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_CMUX = CLBLL_L_X102Y121_SLICE_X161Y121_C5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A = CLBLL_L_X102Y122_SLICE_X160Y122_AO6;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B = CLBLL_L_X102Y122_SLICE_X160Y122_BO6;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C = CLBLL_L_X102Y122_SLICE_X160Y122_CO6;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D = CLBLL_L_X102Y122_SLICE_X160Y122_DO6;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_AMUX = CLBLL_L_X102Y122_SLICE_X160Y122_A5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_BMUX = CLBLL_L_X102Y122_SLICE_X160Y122_B5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_CMUX = CLBLL_L_X102Y122_SLICE_X160Y122_C5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A = CLBLL_L_X102Y122_SLICE_X161Y122_AO6;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B = CLBLL_L_X102Y122_SLICE_X161Y122_BO6;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C = CLBLL_L_X102Y122_SLICE_X161Y122_CO6;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D = CLBLL_L_X102Y122_SLICE_X161Y122_DO6;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_AMUX = CLBLL_L_X102Y122_SLICE_X161Y122_A5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_BMUX = CLBLL_L_X102Y122_SLICE_X161Y122_B5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_CMUX = CLBLL_L_X102Y122_SLICE_X161Y122_C5Q;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A = CLBLL_L_X102Y123_SLICE_X160Y123_AO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B = CLBLL_L_X102Y123_SLICE_X160Y123_BO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C = CLBLL_L_X102Y123_SLICE_X160Y123_CO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D = CLBLL_L_X102Y123_SLICE_X160Y123_DO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_BMUX = CLBLL_L_X102Y123_SLICE_X160Y123_B5Q;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A = CLBLL_L_X102Y123_SLICE_X161Y123_AO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B = CLBLL_L_X102Y123_SLICE_X161Y123_BO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C = CLBLL_L_X102Y123_SLICE_X161Y123_CO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D = CLBLL_L_X102Y123_SLICE_X161Y123_DO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_AMUX = CLBLL_L_X102Y123_SLICE_X161Y123_A5Q;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_DMUX = CLBLL_L_X102Y123_SLICE_X161Y123_DO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A = CLBLL_L_X102Y124_SLICE_X160Y124_AO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B = CLBLL_L_X102Y124_SLICE_X160Y124_BO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C = CLBLL_L_X102Y124_SLICE_X160Y124_CO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D = CLBLL_L_X102Y124_SLICE_X160Y124_DO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_AMUX = CLBLL_L_X102Y124_SLICE_X160Y124_A5Q;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_CMUX = CLBLL_L_X102Y124_SLICE_X160Y124_C5Q;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_DMUX = CLBLL_L_X102Y124_SLICE_X160Y124_D5Q;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A = CLBLL_L_X102Y124_SLICE_X161Y124_AO6;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B = CLBLL_L_X102Y124_SLICE_X161Y124_BO6;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C = CLBLL_L_X102Y124_SLICE_X161Y124_CO6;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D = CLBLL_L_X102Y124_SLICE_X161Y124_DO6;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_AMUX = CLBLL_L_X102Y124_SLICE_X161Y124_A5Q;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_BMUX = CLBLL_L_X102Y124_SLICE_X161Y124_B5Q;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A = CLBLL_L_X102Y125_SLICE_X160Y125_AO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B = CLBLL_L_X102Y125_SLICE_X160Y125_BO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C = CLBLL_L_X102Y125_SLICE_X160Y125_CO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D = CLBLL_L_X102Y125_SLICE_X160Y125_DO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_BMUX = CLBLL_L_X102Y125_SLICE_X160Y125_B5Q;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A = CLBLL_L_X102Y125_SLICE_X161Y125_AO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B = CLBLL_L_X102Y125_SLICE_X161Y125_BO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C = CLBLL_L_X102Y125_SLICE_X161Y125_CO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D = CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_BMUX = CLBLL_L_X102Y125_SLICE_X161Y125_B5Q;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_CMUX = CLBLL_L_X102Y125_SLICE_X161Y125_C5Q;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_DMUX = CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A = CLBLL_L_X102Y126_SLICE_X160Y126_AO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B = CLBLL_L_X102Y126_SLICE_X160Y126_BO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C = CLBLL_L_X102Y126_SLICE_X160Y126_CO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D = CLBLL_L_X102Y126_SLICE_X160Y126_DO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_AMUX = CLBLL_L_X102Y126_SLICE_X160Y126_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_CMUX = CLBLL_L_X102Y126_SLICE_X160Y126_C5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A = CLBLL_L_X102Y126_SLICE_X161Y126_AO6;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B = CLBLL_L_X102Y126_SLICE_X161Y126_BO6;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C = CLBLL_L_X102Y126_SLICE_X161Y126_CO6;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D = CLBLL_L_X102Y126_SLICE_X161Y126_DO6;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_AMUX = CLBLL_L_X102Y126_SLICE_X161Y126_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_BMUX = CLBLL_L_X102Y126_SLICE_X161Y126_B5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_CMUX = CLBLL_L_X102Y126_SLICE_X161Y126_C5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_DMUX = CLBLL_L_X102Y126_SLICE_X161Y126_D5Q;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A = CLBLL_L_X102Y127_SLICE_X160Y127_AO6;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B = CLBLL_L_X102Y127_SLICE_X160Y127_BO6;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C = CLBLL_L_X102Y127_SLICE_X160Y127_CO6;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D = CLBLL_L_X102Y127_SLICE_X160Y127_DO6;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_AMUX = CLBLL_L_X102Y127_SLICE_X160Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_CMUX = CLBLL_L_X102Y127_SLICE_X160Y127_C5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A = CLBLL_L_X102Y127_SLICE_X161Y127_AO6;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B = CLBLL_L_X102Y127_SLICE_X161Y127_BO6;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C = CLBLL_L_X102Y127_SLICE_X161Y127_CO6;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D = CLBLL_L_X102Y127_SLICE_X161Y127_DO6;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_AMUX = CLBLL_L_X102Y127_SLICE_X161Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_BMUX = CLBLL_L_X102Y127_SLICE_X161Y127_B5Q;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A = CLBLL_L_X102Y128_SLICE_X160Y128_AO6;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B = CLBLL_L_X102Y128_SLICE_X160Y128_BO6;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C = CLBLL_L_X102Y128_SLICE_X160Y128_CO6;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D = CLBLL_L_X102Y128_SLICE_X160Y128_DO6;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A = CLBLL_L_X102Y128_SLICE_X161Y128_AO6;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B = CLBLL_L_X102Y128_SLICE_X161Y128_BO6;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C = CLBLL_L_X102Y128_SLICE_X161Y128_CO6;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D = CLBLL_L_X102Y128_SLICE_X161Y128_DO6;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_BMUX = CLBLL_L_X102Y128_SLICE_X161Y128_B5Q;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A = CLBLL_L_X102Y129_SLICE_X160Y129_AO6;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B = CLBLL_L_X102Y129_SLICE_X160Y129_BO6;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C = CLBLL_L_X102Y129_SLICE_X160Y129_CO6;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D = CLBLL_L_X102Y129_SLICE_X160Y129_DO6;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_AMUX = CLBLL_L_X102Y129_SLICE_X160Y129_A5Q;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_CMUX = CLBLL_L_X102Y129_SLICE_X160Y129_C5Q;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A = CLBLL_L_X102Y129_SLICE_X161Y129_AO6;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B = CLBLL_L_X102Y129_SLICE_X161Y129_BO6;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C = CLBLL_L_X102Y129_SLICE_X161Y129_CO6;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D = CLBLL_L_X102Y129_SLICE_X161Y129_DO6;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A = CLBLL_L_X102Y130_SLICE_X160Y130_AO6;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B = CLBLL_L_X102Y130_SLICE_X160Y130_BO6;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C = CLBLL_L_X102Y130_SLICE_X160Y130_CO6;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D = CLBLL_L_X102Y130_SLICE_X160Y130_DO6;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_AMUX = CLBLL_L_X102Y130_SLICE_X160Y130_A5Q;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_BMUX = CLBLL_L_X102Y130_SLICE_X160Y130_B5Q;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_CMUX = CLBLL_L_X102Y130_SLICE_X160Y130_CO6;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A = CLBLL_L_X102Y130_SLICE_X161Y130_AO6;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B = CLBLL_L_X102Y130_SLICE_X161Y130_BO6;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C = CLBLL_L_X102Y130_SLICE_X161Y130_CO6;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D = CLBLL_L_X102Y130_SLICE_X161Y130_DO6;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_AMUX = CLBLL_L_X102Y130_SLICE_X161Y130_A5Q;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A = CLBLL_L_X102Y131_SLICE_X160Y131_AO6;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B = CLBLL_L_X102Y131_SLICE_X160Y131_BO6;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C = CLBLL_L_X102Y131_SLICE_X160Y131_CO6;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D = CLBLL_L_X102Y131_SLICE_X160Y131_DO6;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_BMUX = CLBLL_L_X102Y131_SLICE_X160Y131_B5Q;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A = CLBLL_L_X102Y131_SLICE_X161Y131_AO6;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B = CLBLL_L_X102Y131_SLICE_X161Y131_BO6;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C = CLBLL_L_X102Y131_SLICE_X161Y131_CO6;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D = CLBLL_L_X102Y131_SLICE_X161Y131_DO6;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A = CLBLL_L_X102Y134_SLICE_X160Y134_AO6;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B = CLBLL_L_X102Y134_SLICE_X160Y134_BO6;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C = CLBLL_L_X102Y134_SLICE_X160Y134_CO6;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D = CLBLL_L_X102Y134_SLICE_X160Y134_DO6;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_AMUX = CLBLL_L_X102Y134_SLICE_X160Y134_A5Q;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A = CLBLL_L_X102Y134_SLICE_X161Y134_AO6;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B = CLBLL_L_X102Y134_SLICE_X161Y134_BO6;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C = CLBLL_L_X102Y134_SLICE_X161Y134_CO6;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D = CLBLL_L_X102Y134_SLICE_X161Y134_DO6;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A = CLBLL_L_X102Y135_SLICE_X160Y135_AO6;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B = CLBLL_L_X102Y135_SLICE_X160Y135_BO6;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C = CLBLL_L_X102Y135_SLICE_X160Y135_CO6;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D = CLBLL_L_X102Y135_SLICE_X160Y135_DO6;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A = CLBLL_L_X102Y135_SLICE_X161Y135_AO6;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B = CLBLL_L_X102Y135_SLICE_X161Y135_BO6;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C = CLBLL_L_X102Y135_SLICE_X161Y135_CO6;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D = CLBLL_L_X102Y135_SLICE_X161Y135_DO6;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A = CLBLL_L_X102Y136_SLICE_X160Y136_AO6;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B = CLBLL_L_X102Y136_SLICE_X160Y136_BO6;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C = CLBLL_L_X102Y136_SLICE_X160Y136_CO6;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D = CLBLL_L_X102Y136_SLICE_X160Y136_DO6;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_BMUX = CLBLL_L_X102Y136_SLICE_X160Y136_B5Q;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A = CLBLL_L_X102Y136_SLICE_X161Y136_AO6;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B = CLBLL_L_X102Y136_SLICE_X161Y136_BO6;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C = CLBLL_L_X102Y136_SLICE_X161Y136_CO6;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D = CLBLL_L_X102Y136_SLICE_X161Y136_DO6;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A = CLBLL_R_X87Y118_SLICE_X138Y118_AO6;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B = CLBLL_R_X87Y118_SLICE_X138Y118_BO6;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C = CLBLL_R_X87Y118_SLICE_X138Y118_CO6;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D = CLBLL_R_X87Y118_SLICE_X138Y118_DO6;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_BMUX = CLBLL_R_X87Y118_SLICE_X138Y118_B5Q;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A = CLBLL_R_X87Y118_SLICE_X139Y118_AO6;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B = CLBLL_R_X87Y118_SLICE_X139Y118_BO6;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C = CLBLL_R_X87Y118_SLICE_X139Y118_CO6;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D = CLBLL_R_X87Y118_SLICE_X139Y118_DO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A = CLBLM_L_X90Y113_SLICE_X142Y113_AO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B = CLBLM_L_X90Y113_SLICE_X142Y113_BO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C = CLBLM_L_X90Y113_SLICE_X142Y113_CO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D = CLBLM_L_X90Y113_SLICE_X142Y113_DO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_AMUX = CLBLM_L_X90Y113_SLICE_X142Y113_A5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A = CLBLM_L_X90Y113_SLICE_X143Y113_AO6;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B = CLBLM_L_X90Y113_SLICE_X143Y113_BO6;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C = CLBLM_L_X90Y113_SLICE_X143Y113_CO6;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D = CLBLM_L_X90Y113_SLICE_X143Y113_DO6;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_AMUX = CLBLM_L_X90Y113_SLICE_X143Y113_A5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_BMUX = CLBLM_L_X90Y113_SLICE_X143Y113_B5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_CMUX = CLBLM_L_X90Y113_SLICE_X143Y113_C5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A = CLBLM_L_X90Y114_SLICE_X142Y114_AO6;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B = CLBLM_L_X90Y114_SLICE_X142Y114_BO6;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C = CLBLM_L_X90Y114_SLICE_X142Y114_CO6;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D = CLBLM_L_X90Y114_SLICE_X142Y114_DO6;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_AMUX = CLBLM_L_X90Y114_SLICE_X142Y114_A5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_BMUX = CLBLM_L_X90Y114_SLICE_X142Y114_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_CMUX = CLBLM_L_X90Y114_SLICE_X142Y114_C5Q;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A = CLBLM_L_X90Y114_SLICE_X143Y114_AO6;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B = CLBLM_L_X90Y114_SLICE_X143Y114_BO6;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C = CLBLM_L_X90Y114_SLICE_X143Y114_CO6;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D = CLBLM_L_X90Y114_SLICE_X143Y114_DO6;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_AMUX = CLBLM_L_X90Y114_SLICE_X143Y114_A5Q;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_BMUX = CLBLM_L_X90Y114_SLICE_X143Y114_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_CMUX = CLBLM_L_X90Y114_SLICE_X143Y114_CO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A = CLBLM_L_X90Y115_SLICE_X142Y115_AO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B = CLBLM_L_X90Y115_SLICE_X142Y115_BO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C = CLBLM_L_X90Y115_SLICE_X142Y115_CO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D = CLBLM_L_X90Y115_SLICE_X142Y115_DO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_AMUX = CLBLM_L_X90Y115_SLICE_X142Y115_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A = CLBLM_L_X90Y115_SLICE_X143Y115_AO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B = CLBLM_L_X90Y115_SLICE_X143Y115_BO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C = CLBLM_L_X90Y115_SLICE_X143Y115_CO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D = CLBLM_L_X90Y115_SLICE_X143Y115_DO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_AMUX = CLBLM_L_X90Y115_SLICE_X143Y115_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_BMUX = CLBLM_L_X90Y115_SLICE_X143Y115_B5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_CMUX = CLBLM_L_X90Y115_SLICE_X143Y115_C5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_DMUX = CLBLM_L_X90Y115_SLICE_X143Y115_DO6;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A = CLBLM_L_X90Y116_SLICE_X142Y116_AO6;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B = CLBLM_L_X90Y116_SLICE_X142Y116_BO6;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C = CLBLM_L_X90Y116_SLICE_X142Y116_CO6;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D = CLBLM_L_X90Y116_SLICE_X142Y116_DO6;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_AMUX = CLBLM_L_X90Y116_SLICE_X142Y116_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_CMUX = CLBLM_L_X90Y116_SLICE_X142Y116_C5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A = CLBLM_L_X90Y116_SLICE_X143Y116_AO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B = CLBLM_L_X90Y116_SLICE_X143Y116_BO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C = CLBLM_L_X90Y116_SLICE_X143Y116_CO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D = CLBLM_L_X90Y116_SLICE_X143Y116_DO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_AMUX = CLBLM_L_X90Y116_SLICE_X143Y116_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_BMUX = CLBLM_L_X90Y116_SLICE_X143Y116_B5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_CMUX = CLBLM_L_X90Y116_SLICE_X143Y116_C5Q;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A = CLBLM_L_X90Y117_SLICE_X142Y117_AO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B = CLBLM_L_X90Y117_SLICE_X142Y117_BO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C = CLBLM_L_X90Y117_SLICE_X142Y117_CO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D = CLBLM_L_X90Y117_SLICE_X142Y117_DO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_AMUX = CLBLM_L_X90Y117_SLICE_X142Y117_A5Q;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_BMUX = CLBLM_L_X90Y117_SLICE_X142Y117_BO5;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_CMUX = CLBLM_L_X90Y117_SLICE_X142Y117_C5Q;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A = CLBLM_L_X90Y117_SLICE_X143Y117_AO6;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B = CLBLM_L_X90Y117_SLICE_X143Y117_BO6;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C = CLBLM_L_X90Y117_SLICE_X143Y117_CO6;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D = CLBLM_L_X90Y117_SLICE_X143Y117_DO6;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_AMUX = CLBLM_L_X90Y117_SLICE_X143Y117_A5Q;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_BMUX = CLBLM_L_X90Y117_SLICE_X143Y117_B5Q;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A = CLBLM_L_X90Y118_SLICE_X142Y118_AO6;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B = CLBLM_L_X90Y118_SLICE_X142Y118_BO6;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C = CLBLM_L_X90Y118_SLICE_X142Y118_CO6;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D = CLBLM_L_X90Y118_SLICE_X142Y118_DO6;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_AMUX = CLBLM_L_X90Y118_SLICE_X142Y118_A5Q;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_BMUX = CLBLM_L_X90Y118_SLICE_X142Y118_B5Q;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_DMUX = CLBLM_L_X90Y118_SLICE_X142Y118_DO6;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A = CLBLM_L_X90Y118_SLICE_X143Y118_AO6;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B = CLBLM_L_X90Y118_SLICE_X143Y118_BO6;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C = CLBLM_L_X90Y118_SLICE_X143Y118_CO6;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D = CLBLM_L_X90Y118_SLICE_X143Y118_DO6;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_AMUX = CLBLM_L_X90Y118_SLICE_X143Y118_A5Q;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_BMUX = CLBLM_L_X90Y118_SLICE_X143Y118_B5Q;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_DMUX = CLBLM_L_X90Y118_SLICE_X143Y118_DO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A = CLBLM_L_X90Y119_SLICE_X142Y119_AO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B = CLBLM_L_X90Y119_SLICE_X142Y119_BO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C = CLBLM_L_X90Y119_SLICE_X142Y119_CO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D = CLBLM_L_X90Y119_SLICE_X142Y119_DO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_AMUX = CLBLM_L_X90Y119_SLICE_X142Y119_AO5;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_BMUX = CLBLM_L_X90Y119_SLICE_X142Y119_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_CMUX = CLBLM_L_X90Y119_SLICE_X142Y119_C5Q;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A = CLBLM_L_X90Y119_SLICE_X143Y119_AO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B = CLBLM_L_X90Y119_SLICE_X143Y119_BO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C = CLBLM_L_X90Y119_SLICE_X143Y119_CO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D = CLBLM_L_X90Y119_SLICE_X143Y119_DO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_AMUX = CLBLM_L_X90Y119_SLICE_X143Y119_AO5;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_BMUX = CLBLM_L_X90Y119_SLICE_X143Y119_B5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A = CLBLM_L_X90Y120_SLICE_X142Y120_AO6;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B = CLBLM_L_X90Y120_SLICE_X142Y120_BO6;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C = CLBLM_L_X90Y120_SLICE_X142Y120_CO6;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D = CLBLM_L_X90Y120_SLICE_X142Y120_DO6;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_AMUX = CLBLM_L_X90Y120_SLICE_X142Y120_A5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_BMUX = CLBLM_L_X90Y120_SLICE_X142Y120_B5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_CMUX = CLBLM_L_X90Y120_SLICE_X142Y120_CO5;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A = CLBLM_L_X90Y120_SLICE_X143Y120_AO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B = CLBLM_L_X90Y120_SLICE_X143Y120_BO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C = CLBLM_L_X90Y120_SLICE_X143Y120_CO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D = CLBLM_L_X90Y120_SLICE_X143Y120_DO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_AMUX = CLBLM_L_X90Y120_SLICE_X143Y120_A5Q;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_CMUX = CLBLM_L_X90Y120_SLICE_X143Y120_C5Q;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A = CLBLM_L_X90Y121_SLICE_X142Y121_AO6;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B = CLBLM_L_X90Y121_SLICE_X142Y121_BO6;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C = CLBLM_L_X90Y121_SLICE_X142Y121_CO6;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D = CLBLM_L_X90Y121_SLICE_X142Y121_DO6;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_AMUX = CLBLM_L_X90Y121_SLICE_X142Y121_A5Q;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A = CLBLM_L_X90Y121_SLICE_X143Y121_AO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B = CLBLM_L_X90Y121_SLICE_X143Y121_BO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C = CLBLM_L_X90Y121_SLICE_X143Y121_CO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D = CLBLM_L_X90Y121_SLICE_X143Y121_DO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_AMUX = CLBLM_L_X90Y121_SLICE_X143Y121_A5Q;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_BMUX = CLBLM_L_X90Y121_SLICE_X143Y121_BO5;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_CMUX = CLBLM_L_X90Y121_SLICE_X143Y121_C5Q;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A = CLBLM_L_X90Y122_SLICE_X142Y122_AO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B = CLBLM_L_X90Y122_SLICE_X142Y122_BO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C = CLBLM_L_X90Y122_SLICE_X142Y122_CO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D = CLBLM_L_X90Y122_SLICE_X142Y122_DO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_AMUX = CLBLM_L_X90Y122_SLICE_X142Y122_A5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A = CLBLM_L_X90Y122_SLICE_X143Y122_AO6;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B = CLBLM_L_X90Y122_SLICE_X143Y122_BO6;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C = CLBLM_L_X90Y122_SLICE_X143Y122_CO6;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D = CLBLM_L_X90Y122_SLICE_X143Y122_DO6;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_AMUX = CLBLM_L_X90Y122_SLICE_X143Y122_A5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_BMUX = CLBLM_L_X90Y122_SLICE_X143Y122_BO5;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_CMUX = CLBLM_L_X90Y122_SLICE_X143Y122_C5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A = CLBLM_L_X90Y123_SLICE_X142Y123_AO6;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B = CLBLM_L_X90Y123_SLICE_X142Y123_BO6;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C = CLBLM_L_X90Y123_SLICE_X142Y123_CO6;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D = CLBLM_L_X90Y123_SLICE_X142Y123_DO6;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_AMUX = CLBLM_L_X90Y123_SLICE_X142Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_BMUX = CLBLM_L_X90Y123_SLICE_X142Y123_B5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_CMUX = CLBLM_L_X90Y123_SLICE_X142Y123_C5Q;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A = CLBLM_L_X90Y123_SLICE_X143Y123_AO6;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B = CLBLM_L_X90Y123_SLICE_X143Y123_BO6;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C = CLBLM_L_X90Y123_SLICE_X143Y123_CO6;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D = CLBLM_L_X90Y123_SLICE_X143Y123_DO6;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_AMUX = CLBLM_L_X90Y123_SLICE_X143Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_BMUX = CLBLM_L_X90Y123_SLICE_X143Y123_BO5;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_CMUX = CLBLM_L_X90Y123_SLICE_X143Y123_C5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A = CLBLM_L_X90Y124_SLICE_X142Y124_AO6;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B = CLBLM_L_X90Y124_SLICE_X142Y124_BO6;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C = CLBLM_L_X90Y124_SLICE_X142Y124_CO6;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D = CLBLM_L_X90Y124_SLICE_X142Y124_DO6;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_AMUX = CLBLM_L_X90Y124_SLICE_X142Y124_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_BMUX = CLBLM_L_X90Y124_SLICE_X142Y124_BO5;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_CMUX = CLBLM_L_X90Y124_SLICE_X142Y124_C5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A = CLBLM_L_X90Y124_SLICE_X143Y124_AO6;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B = CLBLM_L_X90Y124_SLICE_X143Y124_BO6;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C = CLBLM_L_X90Y124_SLICE_X143Y124_CO6;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D = CLBLM_L_X90Y124_SLICE_X143Y124_DO6;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_BMUX = CLBLM_L_X90Y124_SLICE_X143Y124_B5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_CMUX = CLBLM_L_X90Y124_SLICE_X143Y124_C5Q;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A = CLBLM_L_X90Y125_SLICE_X142Y125_AO6;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B = CLBLM_L_X90Y125_SLICE_X142Y125_BO6;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C = CLBLM_L_X90Y125_SLICE_X142Y125_CO6;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D = CLBLM_L_X90Y125_SLICE_X142Y125_DO6;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_AMUX = CLBLM_L_X90Y125_SLICE_X142Y125_A5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A = CLBLM_L_X90Y125_SLICE_X143Y125_AO6;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B = CLBLM_L_X90Y125_SLICE_X143Y125_BO6;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C = CLBLM_L_X90Y125_SLICE_X143Y125_CO6;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D = CLBLM_L_X90Y125_SLICE_X143Y125_DO6;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_AMUX = CLBLM_L_X90Y125_SLICE_X143Y125_A5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_BMUX = CLBLM_L_X90Y125_SLICE_X143Y125_B5Q;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A = CLBLM_L_X90Y126_SLICE_X142Y126_AO6;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B = CLBLM_L_X90Y126_SLICE_X142Y126_BO6;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C = CLBLM_L_X90Y126_SLICE_X142Y126_CO6;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D = CLBLM_L_X90Y126_SLICE_X142Y126_DO6;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_BMUX = CLBLM_L_X90Y126_SLICE_X142Y126_B5Q;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_CMUX = CLBLM_L_X90Y126_SLICE_X142Y126_C5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A = CLBLM_L_X90Y126_SLICE_X143Y126_AO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B = CLBLM_L_X90Y126_SLICE_X143Y126_BO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C = CLBLM_L_X90Y126_SLICE_X143Y126_CO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D = CLBLM_L_X90Y126_SLICE_X143Y126_DO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_AMUX = CLBLM_L_X90Y126_SLICE_X143Y126_A5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_BMUX = CLBLM_L_X90Y126_SLICE_X143Y126_BO5;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_CMUX = CLBLM_L_X90Y126_SLICE_X143Y126_C5Q;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A = CLBLM_L_X90Y128_SLICE_X142Y128_AO6;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B = CLBLM_L_X90Y128_SLICE_X142Y128_BO6;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C = CLBLM_L_X90Y128_SLICE_X142Y128_CO6;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D = CLBLM_L_X90Y128_SLICE_X142Y128_DO6;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_AMUX = CLBLM_L_X90Y128_SLICE_X142Y128_AO6;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_BMUX = CLBLM_L_X90Y128_SLICE_X142Y128_B5Q;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A = CLBLM_L_X90Y128_SLICE_X143Y128_AO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B = CLBLM_L_X90Y128_SLICE_X143Y128_BO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C = CLBLM_L_X90Y128_SLICE_X143Y128_CO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D = CLBLM_L_X90Y128_SLICE_X143Y128_DO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_AMUX = CLBLM_L_X90Y128_SLICE_X143Y128_A5Q;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_DMUX = CLBLM_L_X90Y128_SLICE_X143Y128_D5Q;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A = CLBLM_L_X90Y129_SLICE_X142Y129_AO6;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B = CLBLM_L_X90Y129_SLICE_X142Y129_BO6;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C = CLBLM_L_X90Y129_SLICE_X142Y129_CO6;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D = CLBLM_L_X90Y129_SLICE_X142Y129_DO6;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_AMUX = CLBLM_L_X90Y129_SLICE_X142Y129_A5Q;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_BMUX = CLBLM_L_X90Y129_SLICE_X142Y129_BO5;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_CMUX = CLBLM_L_X90Y129_SLICE_X142Y129_C5Q;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A = CLBLM_L_X90Y129_SLICE_X143Y129_AO6;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B = CLBLM_L_X90Y129_SLICE_X143Y129_BO6;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C = CLBLM_L_X90Y129_SLICE_X143Y129_CO6;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D = CLBLM_L_X90Y129_SLICE_X143Y129_DO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A = CLBLM_L_X90Y130_SLICE_X142Y130_AO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B = CLBLM_L_X90Y130_SLICE_X142Y130_BO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C = CLBLM_L_X90Y130_SLICE_X142Y130_CO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D = CLBLM_L_X90Y130_SLICE_X142Y130_DO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_AMUX = CLBLM_L_X90Y130_SLICE_X142Y130_A5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_BMUX = CLBLM_L_X90Y130_SLICE_X142Y130_B5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_CMUX = CLBLM_L_X90Y130_SLICE_X142Y130_CO5;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A = CLBLM_L_X90Y130_SLICE_X143Y130_AO6;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B = CLBLM_L_X90Y130_SLICE_X143Y130_BO6;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C = CLBLM_L_X90Y130_SLICE_X143Y130_CO6;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D = CLBLM_L_X90Y130_SLICE_X143Y130_DO6;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A = CLBLM_L_X90Y131_SLICE_X142Y131_AO6;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B = CLBLM_L_X90Y131_SLICE_X142Y131_BO6;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C = CLBLM_L_X90Y131_SLICE_X142Y131_CO6;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D = CLBLM_L_X90Y131_SLICE_X142Y131_DO6;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_AMUX = CLBLM_L_X90Y131_SLICE_X142Y131_A5Q;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_BMUX = CLBLM_L_X90Y131_SLICE_X142Y131_BO5;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_CMUX = CLBLM_L_X90Y131_SLICE_X142Y131_C5Q;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A = CLBLM_L_X90Y131_SLICE_X143Y131_AO6;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B = CLBLM_L_X90Y131_SLICE_X143Y131_BO6;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C = CLBLM_L_X90Y131_SLICE_X143Y131_CO6;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D = CLBLM_L_X90Y131_SLICE_X143Y131_DO6;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A = CLBLM_L_X92Y112_SLICE_X144Y112_AO6;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B = CLBLM_L_X92Y112_SLICE_X144Y112_BO6;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C = CLBLM_L_X92Y112_SLICE_X144Y112_CO6;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D = CLBLM_L_X92Y112_SLICE_X144Y112_DO6;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A = CLBLM_L_X92Y112_SLICE_X145Y112_AO6;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B = CLBLM_L_X92Y112_SLICE_X145Y112_BO6;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C = CLBLM_L_X92Y112_SLICE_X145Y112_CO6;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D = CLBLM_L_X92Y112_SLICE_X145Y112_DO6;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_AMUX = CLBLM_L_X92Y112_SLICE_X145Y112_A5Q;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_BMUX = CLBLM_L_X92Y112_SLICE_X145Y112_B5Q;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A = CLBLM_L_X92Y113_SLICE_X144Y113_AO6;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B = CLBLM_L_X92Y113_SLICE_X144Y113_BO6;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C = CLBLM_L_X92Y113_SLICE_X144Y113_CO6;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D = CLBLM_L_X92Y113_SLICE_X144Y113_DO6;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_AMUX = CLBLM_L_X92Y113_SLICE_X144Y113_A5Q;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_BMUX = CLBLM_L_X92Y113_SLICE_X144Y113_B5Q;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A = CLBLM_L_X92Y113_SLICE_X145Y113_AO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B = CLBLM_L_X92Y113_SLICE_X145Y113_BO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C = CLBLM_L_X92Y113_SLICE_X145Y113_CO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D = CLBLM_L_X92Y113_SLICE_X145Y113_DO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_AMUX = CLBLM_L_X92Y113_SLICE_X145Y113_A5Q;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_BMUX = CLBLM_L_X92Y113_SLICE_X145Y113_B5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A = CLBLM_L_X92Y114_SLICE_X144Y114_AO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B = CLBLM_L_X92Y114_SLICE_X144Y114_BO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C = CLBLM_L_X92Y114_SLICE_X144Y114_CO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D = CLBLM_L_X92Y114_SLICE_X144Y114_DO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_AMUX = CLBLM_L_X92Y114_SLICE_X144Y114_A5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_BMUX = CLBLM_L_X92Y114_SLICE_X144Y114_B5Q;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A = CLBLM_L_X92Y114_SLICE_X145Y114_AO6;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B = CLBLM_L_X92Y114_SLICE_X145Y114_BO6;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C = CLBLM_L_X92Y114_SLICE_X145Y114_CO6;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D = CLBLM_L_X92Y114_SLICE_X145Y114_DO6;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_AMUX = CLBLM_L_X92Y114_SLICE_X145Y114_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A = CLBLM_L_X92Y115_SLICE_X144Y115_AO6;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B = CLBLM_L_X92Y115_SLICE_X144Y115_BO6;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C = CLBLM_L_X92Y115_SLICE_X144Y115_CO6;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D = CLBLM_L_X92Y115_SLICE_X144Y115_DO6;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A = CLBLM_L_X92Y115_SLICE_X145Y115_AO6;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B = CLBLM_L_X92Y115_SLICE_X145Y115_BO6;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C = CLBLM_L_X92Y115_SLICE_X145Y115_CO6;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D = CLBLM_L_X92Y115_SLICE_X145Y115_DO6;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_AMUX = CLBLM_L_X92Y115_SLICE_X145Y115_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_BMUX = CLBLM_L_X92Y115_SLICE_X145Y115_B5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A = CLBLM_L_X92Y116_SLICE_X144Y116_AO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B = CLBLM_L_X92Y116_SLICE_X144Y116_BO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C = CLBLM_L_X92Y116_SLICE_X144Y116_CO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D = CLBLM_L_X92Y116_SLICE_X144Y116_DO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_AMUX = CLBLM_L_X92Y116_SLICE_X144Y116_A5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_BMUX = CLBLM_L_X92Y116_SLICE_X144Y116_B5Q;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A = CLBLM_L_X92Y116_SLICE_X145Y116_AO6;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B = CLBLM_L_X92Y116_SLICE_X145Y116_BO6;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C = CLBLM_L_X92Y116_SLICE_X145Y116_CO6;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D = CLBLM_L_X92Y116_SLICE_X145Y116_DO6;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_AMUX = CLBLM_L_X92Y116_SLICE_X145Y116_A5Q;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_BMUX = CLBLM_L_X92Y116_SLICE_X145Y116_B5Q;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A = CLBLM_L_X92Y118_SLICE_X144Y118_AO6;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B = CLBLM_L_X92Y118_SLICE_X144Y118_BO6;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C = CLBLM_L_X92Y118_SLICE_X144Y118_CO6;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D = CLBLM_L_X92Y118_SLICE_X144Y118_DO6;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_AMUX = CLBLM_L_X92Y118_SLICE_X144Y118_A5Q;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A = CLBLM_L_X92Y118_SLICE_X145Y118_AO6;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B = CLBLM_L_X92Y118_SLICE_X145Y118_BO6;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C = CLBLM_L_X92Y118_SLICE_X145Y118_CO6;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D = CLBLM_L_X92Y118_SLICE_X145Y118_DO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A = CLBLM_L_X92Y119_SLICE_X144Y119_AO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B = CLBLM_L_X92Y119_SLICE_X144Y119_BO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C = CLBLM_L_X92Y119_SLICE_X144Y119_CO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D = CLBLM_L_X92Y119_SLICE_X144Y119_DO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_AMUX = CLBLM_L_X92Y119_SLICE_X144Y119_A5Q;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_BMUX = CLBLM_L_X92Y119_SLICE_X144Y119_BO5;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_CMUX = CLBLM_L_X92Y119_SLICE_X144Y119_C5Q;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A = CLBLM_L_X92Y119_SLICE_X145Y119_AO6;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B = CLBLM_L_X92Y119_SLICE_X145Y119_BO6;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C = CLBLM_L_X92Y119_SLICE_X145Y119_CO6;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D = CLBLM_L_X92Y119_SLICE_X145Y119_DO6;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_AMUX = CLBLM_L_X92Y119_SLICE_X145Y119_A5Q;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_BMUX = CLBLM_L_X92Y119_SLICE_X145Y119_B5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A = CLBLM_L_X92Y120_SLICE_X144Y120_AO6;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B = CLBLM_L_X92Y120_SLICE_X144Y120_BO6;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C = CLBLM_L_X92Y120_SLICE_X144Y120_CO6;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D = CLBLM_L_X92Y120_SLICE_X144Y120_DO6;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_AMUX = CLBLM_L_X92Y120_SLICE_X144Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_BMUX = CLBLM_L_X92Y120_SLICE_X144Y120_B5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A = CLBLM_L_X92Y120_SLICE_X145Y120_AO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B = CLBLM_L_X92Y120_SLICE_X145Y120_BO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C = CLBLM_L_X92Y120_SLICE_X145Y120_CO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D = CLBLM_L_X92Y120_SLICE_X145Y120_DO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_AMUX = CLBLM_L_X92Y120_SLICE_X145Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_BMUX = CLBLM_L_X92Y120_SLICE_X145Y120_BO5;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_CMUX = CLBLM_L_X92Y120_SLICE_X145Y120_C5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A = CLBLM_L_X92Y121_SLICE_X144Y121_AO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B = CLBLM_L_X92Y121_SLICE_X144Y121_BO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C = CLBLM_L_X92Y121_SLICE_X144Y121_CO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D = CLBLM_L_X92Y121_SLICE_X144Y121_DO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_AMUX = CLBLM_L_X92Y121_SLICE_X144Y121_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_DMUX = CLBLM_L_X92Y121_SLICE_X144Y121_D5Q;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A = CLBLM_L_X92Y121_SLICE_X145Y121_AO6;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B = CLBLM_L_X92Y121_SLICE_X145Y121_BO6;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C = CLBLM_L_X92Y121_SLICE_X145Y121_CO6;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D = CLBLM_L_X92Y121_SLICE_X145Y121_DO6;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_AMUX = CLBLM_L_X92Y121_SLICE_X145Y121_AO6;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_BMUX = CLBLM_L_X92Y121_SLICE_X145Y121_B5Q;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_CMUX = CLBLM_L_X92Y121_SLICE_X145Y121_C5Q;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A = CLBLM_L_X92Y122_SLICE_X144Y122_AO6;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B = CLBLM_L_X92Y122_SLICE_X144Y122_BO6;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C = CLBLM_L_X92Y122_SLICE_X144Y122_CO6;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D = CLBLM_L_X92Y122_SLICE_X144Y122_DO6;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_BMUX = CLBLM_L_X92Y122_SLICE_X144Y122_B5Q;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_CMUX = CLBLM_L_X92Y122_SLICE_X144Y122_C5Q;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A = CLBLM_L_X92Y122_SLICE_X145Y122_AO6;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B = CLBLM_L_X92Y122_SLICE_X145Y122_BO6;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C = CLBLM_L_X92Y122_SLICE_X145Y122_CO6;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D = CLBLM_L_X92Y122_SLICE_X145Y122_DO6;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_BMUX = CLBLM_L_X92Y122_SLICE_X145Y122_B5Q;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_CMUX = CLBLM_L_X92Y122_SLICE_X145Y122_C5Q;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A = CLBLM_L_X92Y123_SLICE_X144Y123_AO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B = CLBLM_L_X92Y123_SLICE_X144Y123_BO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C = CLBLM_L_X92Y123_SLICE_X144Y123_CO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D = CLBLM_L_X92Y123_SLICE_X144Y123_DO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_AMUX = CLBLM_L_X92Y123_SLICE_X144Y123_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_DMUX = CLBLM_L_X92Y123_SLICE_X144Y123_D5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A = CLBLM_L_X92Y123_SLICE_X145Y123_AO6;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B = CLBLM_L_X92Y123_SLICE_X145Y123_BO6;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C = CLBLM_L_X92Y123_SLICE_X145Y123_CO6;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D = CLBLM_L_X92Y123_SLICE_X145Y123_DO6;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_AMUX = CLBLM_L_X92Y123_SLICE_X145Y123_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_BMUX = CLBLM_L_X92Y123_SLICE_X145Y123_B5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_DMUX = CLBLM_L_X92Y123_SLICE_X145Y123_DO5;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A = CLBLM_L_X92Y124_SLICE_X144Y124_AO6;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B = CLBLM_L_X92Y124_SLICE_X144Y124_BO6;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C = CLBLM_L_X92Y124_SLICE_X144Y124_CO6;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D = CLBLM_L_X92Y124_SLICE_X144Y124_DO6;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_AMUX = CLBLM_L_X92Y124_SLICE_X144Y124_A5Q;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_BMUX = CLBLM_L_X92Y124_SLICE_X144Y124_BO5;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_CMUX = CLBLM_L_X92Y124_SLICE_X144Y124_C5Q;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A = CLBLM_L_X92Y124_SLICE_X145Y124_AO6;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B = CLBLM_L_X92Y124_SLICE_X145Y124_BO6;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C = CLBLM_L_X92Y124_SLICE_X145Y124_CO6;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D = CLBLM_L_X92Y124_SLICE_X145Y124_DO6;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_AMUX = CLBLM_L_X92Y124_SLICE_X145Y124_A5Q;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A = CLBLM_L_X92Y125_SLICE_X144Y125_AO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B = CLBLM_L_X92Y125_SLICE_X144Y125_BO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C = CLBLM_L_X92Y125_SLICE_X144Y125_CO6;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D = CLBLM_L_X92Y125_SLICE_X144Y125_DO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A = CLBLM_L_X92Y125_SLICE_X145Y125_AO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B = CLBLM_L_X92Y125_SLICE_X145Y125_BO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C = CLBLM_L_X92Y125_SLICE_X145Y125_CO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D = CLBLM_L_X92Y125_SLICE_X145Y125_DO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_AMUX = CLBLM_L_X92Y125_SLICE_X145Y125_A5Q;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_BMUX = CLBLM_L_X92Y125_SLICE_X145Y125_BO5;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_CMUX = CLBLM_L_X92Y125_SLICE_X145Y125_C5Q;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A = CLBLM_L_X92Y126_SLICE_X144Y126_AO6;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B = CLBLM_L_X92Y126_SLICE_X144Y126_BO6;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C = CLBLM_L_X92Y126_SLICE_X144Y126_CO6;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D = CLBLM_L_X92Y126_SLICE_X144Y126_DO6;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A = CLBLM_L_X92Y126_SLICE_X145Y126_AO6;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B = CLBLM_L_X92Y126_SLICE_X145Y126_BO6;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C = CLBLM_L_X92Y126_SLICE_X145Y126_CO6;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D = CLBLM_L_X92Y126_SLICE_X145Y126_DO6;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_AMUX = CLBLM_L_X92Y126_SLICE_X145Y126_AO5;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_BMUX = CLBLM_L_X92Y126_SLICE_X145Y126_B5Q;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_CMUX = CLBLM_L_X92Y126_SLICE_X145Y126_C5Q;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A = CLBLM_L_X92Y127_SLICE_X144Y127_AO6;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B = CLBLM_L_X92Y127_SLICE_X144Y127_BO6;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C = CLBLM_L_X92Y127_SLICE_X144Y127_CO6;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D = CLBLM_L_X92Y127_SLICE_X144Y127_DO6;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A = CLBLM_L_X92Y127_SLICE_X145Y127_AO6;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B = CLBLM_L_X92Y127_SLICE_X145Y127_BO6;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C = CLBLM_L_X92Y127_SLICE_X145Y127_CO6;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D = CLBLM_L_X92Y127_SLICE_X145Y127_DO6;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_BMUX = CLBLM_L_X92Y127_SLICE_X145Y127_B5Q;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A = CLBLM_L_X92Y128_SLICE_X144Y128_AO6;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B = CLBLM_L_X92Y128_SLICE_X144Y128_BO6;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C = CLBLM_L_X92Y128_SLICE_X144Y128_CO6;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D = CLBLM_L_X92Y128_SLICE_X144Y128_DO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A = CLBLM_L_X92Y128_SLICE_X145Y128_AO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B = CLBLM_L_X92Y128_SLICE_X145Y128_BO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C = CLBLM_L_X92Y128_SLICE_X145Y128_CO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D = CLBLM_L_X92Y128_SLICE_X145Y128_DO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_AMUX = CLBLM_L_X92Y128_SLICE_X145Y128_A5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_BMUX = CLBLM_L_X92Y128_SLICE_X145Y128_BO5;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_CMUX = CLBLM_L_X92Y128_SLICE_X145Y128_C5Q;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A = CLBLM_L_X92Y129_SLICE_X144Y129_AO6;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B = CLBLM_L_X92Y129_SLICE_X144Y129_BO6;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C = CLBLM_L_X92Y129_SLICE_X144Y129_CO6;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D = CLBLM_L_X92Y129_SLICE_X144Y129_DO6;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A = CLBLM_L_X92Y129_SLICE_X145Y129_AO6;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B = CLBLM_L_X92Y129_SLICE_X145Y129_BO6;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C = CLBLM_L_X92Y129_SLICE_X145Y129_CO6;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D = CLBLM_L_X92Y129_SLICE_X145Y129_DO6;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_AMUX = CLBLM_L_X92Y129_SLICE_X145Y129_A5Q;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_BMUX = CLBLM_L_X92Y129_SLICE_X145Y129_BO5;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_CMUX = CLBLM_L_X92Y129_SLICE_X145Y129_C5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A = CLBLM_L_X92Y131_SLICE_X144Y131_AO6;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B = CLBLM_L_X92Y131_SLICE_X144Y131_BO6;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C = CLBLM_L_X92Y131_SLICE_X144Y131_CO6;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D = CLBLM_L_X92Y131_SLICE_X144Y131_DO6;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_AMUX = CLBLM_L_X92Y131_SLICE_X144Y131_A5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_BMUX = CLBLM_L_X92Y131_SLICE_X144Y131_B5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_CMUX = CLBLM_L_X92Y131_SLICE_X144Y131_C5Q;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A = CLBLM_L_X92Y131_SLICE_X145Y131_AO6;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B = CLBLM_L_X92Y131_SLICE_X145Y131_BO6;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C = CLBLM_L_X92Y131_SLICE_X145Y131_CO6;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D = CLBLM_L_X92Y131_SLICE_X145Y131_DO6;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_AMUX = CLBLM_L_X92Y131_SLICE_X145Y131_A5Q;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_BMUX = CLBLM_L_X92Y131_SLICE_X145Y131_BO5;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A = CLBLM_L_X92Y132_SLICE_X144Y132_AO6;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B = CLBLM_L_X92Y132_SLICE_X144Y132_BO6;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C = CLBLM_L_X92Y132_SLICE_X144Y132_CO6;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D = CLBLM_L_X92Y132_SLICE_X144Y132_DO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A = CLBLM_L_X92Y132_SLICE_X145Y132_AO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B = CLBLM_L_X92Y132_SLICE_X145Y132_BO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C = CLBLM_L_X92Y132_SLICE_X145Y132_CO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D = CLBLM_L_X92Y132_SLICE_X145Y132_DO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_AMUX = CLBLM_L_X92Y132_SLICE_X145Y132_A5Q;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_BMUX = CLBLM_L_X92Y132_SLICE_X145Y132_BO5;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_CMUX = CLBLM_L_X92Y132_SLICE_X145Y132_C5Q;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A = CLBLM_L_X94Y111_SLICE_X148Y111_AO6;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B = CLBLM_L_X94Y111_SLICE_X148Y111_BO6;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C = CLBLM_L_X94Y111_SLICE_X148Y111_CO6;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D = CLBLM_L_X94Y111_SLICE_X148Y111_DO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A = CLBLM_L_X94Y111_SLICE_X149Y111_AO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B = CLBLM_L_X94Y111_SLICE_X149Y111_BO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C = CLBLM_L_X94Y111_SLICE_X149Y111_CO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D = CLBLM_L_X94Y111_SLICE_X149Y111_DO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_AMUX = CLBLM_L_X94Y111_SLICE_X149Y111_A5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_BMUX = CLBLM_L_X94Y111_SLICE_X149Y111_B5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_CMUX = CLBLM_L_X94Y111_SLICE_X149Y111_CO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A = CLBLM_L_X94Y112_SLICE_X148Y112_AO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B = CLBLM_L_X94Y112_SLICE_X148Y112_BO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C = CLBLM_L_X94Y112_SLICE_X148Y112_CO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D = CLBLM_L_X94Y112_SLICE_X148Y112_DO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_AMUX = CLBLM_L_X94Y112_SLICE_X148Y112_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_BMUX = CLBLM_L_X94Y112_SLICE_X148Y112_B5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A = CLBLM_L_X94Y112_SLICE_X149Y112_AO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B = CLBLM_L_X94Y112_SLICE_X149Y112_BO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C = CLBLM_L_X94Y112_SLICE_X149Y112_CO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D = CLBLM_L_X94Y112_SLICE_X149Y112_DO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_AMUX = CLBLM_L_X94Y112_SLICE_X149Y112_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_BMUX = CLBLM_L_X94Y112_SLICE_X149Y112_B5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_CMUX = CLBLM_L_X94Y112_SLICE_X149Y112_CO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A = CLBLM_L_X94Y113_SLICE_X148Y113_AO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B = CLBLM_L_X94Y113_SLICE_X148Y113_BO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C = CLBLM_L_X94Y113_SLICE_X148Y113_CO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D = CLBLM_L_X94Y113_SLICE_X148Y113_DO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_AMUX = CLBLM_L_X94Y113_SLICE_X148Y113_A5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_BMUX = CLBLM_L_X94Y113_SLICE_X148Y113_B5Q;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A = CLBLM_L_X94Y113_SLICE_X149Y113_AO6;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B = CLBLM_L_X94Y113_SLICE_X149Y113_BO6;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C = CLBLM_L_X94Y113_SLICE_X149Y113_CO6;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D = CLBLM_L_X94Y113_SLICE_X149Y113_DO6;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_AMUX = CLBLM_L_X94Y113_SLICE_X149Y113_A5Q;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_BMUX = CLBLM_L_X94Y113_SLICE_X149Y113_BO6;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A = CLBLM_L_X94Y114_SLICE_X148Y114_AO6;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B = CLBLM_L_X94Y114_SLICE_X148Y114_BO6;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C = CLBLM_L_X94Y114_SLICE_X148Y114_CO6;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D = CLBLM_L_X94Y114_SLICE_X148Y114_DO6;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_AMUX = CLBLM_L_X94Y114_SLICE_X148Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_BMUX = CLBLM_L_X94Y114_SLICE_X148Y114_B5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A = CLBLM_L_X94Y114_SLICE_X149Y114_AO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B = CLBLM_L_X94Y114_SLICE_X149Y114_BO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C = CLBLM_L_X94Y114_SLICE_X149Y114_CO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D = CLBLM_L_X94Y114_SLICE_X149Y114_DO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_AMUX = CLBLM_L_X94Y114_SLICE_X149Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_BMUX = CLBLM_L_X94Y114_SLICE_X149Y114_B5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_DMUX = CLBLM_L_X94Y114_SLICE_X149Y114_DO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A = CLBLM_L_X94Y115_SLICE_X148Y115_AO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B = CLBLM_L_X94Y115_SLICE_X148Y115_BO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C = CLBLM_L_X94Y115_SLICE_X148Y115_CO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D = CLBLM_L_X94Y115_SLICE_X148Y115_DO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_AMUX = CLBLM_L_X94Y115_SLICE_X148Y115_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_BMUX = CLBLM_L_X94Y115_SLICE_X148Y115_B5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_CMUX = CLBLM_L_X94Y115_SLICE_X148Y115_C5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_DMUX = CLBLM_L_X94Y115_SLICE_X148Y115_DO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A = CLBLM_L_X94Y115_SLICE_X149Y115_AO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B = CLBLM_L_X94Y115_SLICE_X149Y115_BO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C = CLBLM_L_X94Y115_SLICE_X149Y115_CO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D = CLBLM_L_X94Y115_SLICE_X149Y115_DO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_AMUX = CLBLM_L_X94Y115_SLICE_X149Y115_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_BMUX = CLBLM_L_X94Y115_SLICE_X149Y115_B5Q;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A = CLBLM_L_X94Y116_SLICE_X148Y116_AO6;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B = CLBLM_L_X94Y116_SLICE_X148Y116_BO6;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C = CLBLM_L_X94Y116_SLICE_X148Y116_CO6;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D = CLBLM_L_X94Y116_SLICE_X148Y116_DO6;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_AMUX = CLBLM_L_X94Y116_SLICE_X148Y116_A5Q;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_BMUX = CLBLM_L_X94Y116_SLICE_X148Y116_B5Q;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_DMUX = CLBLM_L_X94Y116_SLICE_X148Y116_DO6;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A = CLBLM_L_X94Y116_SLICE_X149Y116_AO6;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B = CLBLM_L_X94Y116_SLICE_X149Y116_BO6;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C = CLBLM_L_X94Y116_SLICE_X149Y116_CO6;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D = CLBLM_L_X94Y116_SLICE_X149Y116_DO6;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_AMUX = CLBLM_L_X94Y116_SLICE_X149Y116_A5Q;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_BMUX = CLBLM_L_X94Y116_SLICE_X149Y116_B5Q;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_CMUX = CLBLM_L_X94Y116_SLICE_X149Y116_C5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A = CLBLM_L_X94Y117_SLICE_X148Y117_AO6;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B = CLBLM_L_X94Y117_SLICE_X148Y117_BO6;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C = CLBLM_L_X94Y117_SLICE_X148Y117_CO6;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D = CLBLM_L_X94Y117_SLICE_X148Y117_DO6;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_AMUX = CLBLM_L_X94Y117_SLICE_X148Y117_A5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_BMUX = CLBLM_L_X94Y117_SLICE_X148Y117_B5Q;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A = CLBLM_L_X94Y117_SLICE_X149Y117_AO6;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B = CLBLM_L_X94Y117_SLICE_X149Y117_BO6;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C = CLBLM_L_X94Y117_SLICE_X149Y117_CO6;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D = CLBLM_L_X94Y117_SLICE_X149Y117_DO6;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_AMUX = CLBLM_L_X94Y117_SLICE_X149Y117_A5Q;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_BMUX = CLBLM_L_X94Y117_SLICE_X149Y117_B5Q;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A = CLBLM_L_X94Y118_SLICE_X148Y118_AO6;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B = CLBLM_L_X94Y118_SLICE_X148Y118_BO6;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C = CLBLM_L_X94Y118_SLICE_X148Y118_CO6;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D = CLBLM_L_X94Y118_SLICE_X148Y118_DO6;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_AMUX = CLBLM_L_X94Y118_SLICE_X148Y118_A5Q;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A = CLBLM_L_X94Y118_SLICE_X149Y118_AO6;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B = CLBLM_L_X94Y118_SLICE_X149Y118_BO6;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C = CLBLM_L_X94Y118_SLICE_X149Y118_CO6;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D = CLBLM_L_X94Y118_SLICE_X149Y118_DO6;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_AMUX = CLBLM_L_X94Y118_SLICE_X149Y118_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A = CLBLM_L_X94Y119_SLICE_X148Y119_AO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B = CLBLM_L_X94Y119_SLICE_X148Y119_BO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C = CLBLM_L_X94Y119_SLICE_X148Y119_CO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D = CLBLM_L_X94Y119_SLICE_X148Y119_DO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_AMUX = CLBLM_L_X94Y119_SLICE_X148Y119_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_CMUX = CLBLM_L_X94Y119_SLICE_X148Y119_CO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A = CLBLM_L_X94Y119_SLICE_X149Y119_AO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B = CLBLM_L_X94Y119_SLICE_X149Y119_BO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C = CLBLM_L_X94Y119_SLICE_X149Y119_CO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D = CLBLM_L_X94Y119_SLICE_X149Y119_DO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_AMUX = CLBLM_L_X94Y119_SLICE_X149Y119_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_BMUX = CLBLM_L_X94Y119_SLICE_X149Y119_B5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A = CLBLM_L_X94Y120_SLICE_X148Y120_AO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B = CLBLM_L_X94Y120_SLICE_X148Y120_BO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C = CLBLM_L_X94Y120_SLICE_X148Y120_CO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D = CLBLM_L_X94Y120_SLICE_X148Y120_DO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_AMUX = CLBLM_L_X94Y120_SLICE_X148Y120_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_BMUX = CLBLM_L_X94Y120_SLICE_X148Y120_B5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_CMUX = CLBLM_L_X94Y120_SLICE_X148Y120_C5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A = CLBLM_L_X94Y120_SLICE_X149Y120_AO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B = CLBLM_L_X94Y120_SLICE_X149Y120_BO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C = CLBLM_L_X94Y120_SLICE_X149Y120_CO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D = CLBLM_L_X94Y120_SLICE_X149Y120_DO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_AMUX = CLBLM_L_X94Y120_SLICE_X149Y120_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_BMUX = CLBLM_L_X94Y120_SLICE_X149Y120_B5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_CMUX = CLBLM_L_X94Y120_SLICE_X149Y120_CO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A = CLBLM_L_X94Y121_SLICE_X148Y121_AO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B = CLBLM_L_X94Y121_SLICE_X148Y121_BO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C = CLBLM_L_X94Y121_SLICE_X148Y121_CO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D = CLBLM_L_X94Y121_SLICE_X148Y121_DO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_AMUX = CLBLM_L_X94Y121_SLICE_X148Y121_A5Q;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_BMUX = CLBLM_L_X94Y121_SLICE_X148Y121_BO5;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_CMUX = CLBLM_L_X94Y121_SLICE_X148Y121_C5Q;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A = CLBLM_L_X94Y121_SLICE_X149Y121_AO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B = CLBLM_L_X94Y121_SLICE_X149Y121_BO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C = CLBLM_L_X94Y121_SLICE_X149Y121_CO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D = CLBLM_L_X94Y121_SLICE_X149Y121_DO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_AMUX = CLBLM_L_X94Y121_SLICE_X149Y121_A5Q;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A = CLBLM_L_X94Y122_SLICE_X148Y122_AO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B = CLBLM_L_X94Y122_SLICE_X148Y122_BO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C = CLBLM_L_X94Y122_SLICE_X148Y122_CO6;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D = CLBLM_L_X94Y122_SLICE_X148Y122_DO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A = CLBLM_L_X94Y122_SLICE_X149Y122_AO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B = CLBLM_L_X94Y122_SLICE_X149Y122_BO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C = CLBLM_L_X94Y122_SLICE_X149Y122_CO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D = CLBLM_L_X94Y122_SLICE_X149Y122_DO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_AMUX = CLBLM_L_X94Y122_SLICE_X149Y122_A5Q;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_BMUX = CLBLM_L_X94Y122_SLICE_X149Y122_B5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A = CLBLM_L_X94Y123_SLICE_X148Y123_AO6;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B = CLBLM_L_X94Y123_SLICE_X148Y123_BO6;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C = CLBLM_L_X94Y123_SLICE_X148Y123_CO6;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D = CLBLM_L_X94Y123_SLICE_X148Y123_DO6;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_AMUX = CLBLM_L_X94Y123_SLICE_X148Y123_A5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_BMUX = CLBLM_L_X94Y123_SLICE_X148Y123_BO5;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_CMUX = CLBLM_L_X94Y123_SLICE_X148Y123_C5Q;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A = CLBLM_L_X94Y123_SLICE_X149Y123_AO6;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B = CLBLM_L_X94Y123_SLICE_X149Y123_BO6;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C = CLBLM_L_X94Y123_SLICE_X149Y123_CO6;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D = CLBLM_L_X94Y123_SLICE_X149Y123_DO6;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A = CLBLM_L_X94Y124_SLICE_X148Y124_AO6;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B = CLBLM_L_X94Y124_SLICE_X148Y124_BO6;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C = CLBLM_L_X94Y124_SLICE_X148Y124_CO6;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D = CLBLM_L_X94Y124_SLICE_X148Y124_DO6;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_AMUX = CLBLM_L_X94Y124_SLICE_X148Y124_A5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_BMUX = CLBLM_L_X94Y124_SLICE_X148Y124_B5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_CMUX = CLBLM_L_X94Y124_SLICE_X148Y124_C5Q;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A = CLBLM_L_X94Y124_SLICE_X149Y124_AO6;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B = CLBLM_L_X94Y124_SLICE_X149Y124_BO6;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C = CLBLM_L_X94Y124_SLICE_X149Y124_CO6;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D = CLBLM_L_X94Y124_SLICE_X149Y124_DO6;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_AMUX = CLBLM_L_X94Y124_SLICE_X149Y124_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A = CLBLM_L_X94Y125_SLICE_X148Y125_AO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B = CLBLM_L_X94Y125_SLICE_X148Y125_BO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C = CLBLM_L_X94Y125_SLICE_X148Y125_CO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D = CLBLM_L_X94Y125_SLICE_X148Y125_DO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_AMUX = CLBLM_L_X94Y125_SLICE_X148Y125_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_BMUX = CLBLM_L_X94Y125_SLICE_X148Y125_B5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_CMUX = CLBLM_L_X94Y125_SLICE_X148Y125_CO6;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A = CLBLM_L_X94Y125_SLICE_X149Y125_AO6;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B = CLBLM_L_X94Y125_SLICE_X149Y125_BO6;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C = CLBLM_L_X94Y125_SLICE_X149Y125_CO6;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D = CLBLM_L_X94Y125_SLICE_X149Y125_DO6;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_AMUX = CLBLM_L_X94Y125_SLICE_X149Y125_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_BMUX = CLBLM_L_X94Y125_SLICE_X149Y125_BO5;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_CMUX = CLBLM_L_X94Y125_SLICE_X149Y125_C5Q;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_DMUX = CLBLM_L_X94Y125_SLICE_X149Y125_D5Q;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A = CLBLM_L_X94Y126_SLICE_X148Y126_AO6;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B = CLBLM_L_X94Y126_SLICE_X148Y126_BO6;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C = CLBLM_L_X94Y126_SLICE_X148Y126_CO6;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D = CLBLM_L_X94Y126_SLICE_X148Y126_DO6;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A = CLBLM_L_X94Y126_SLICE_X149Y126_AO6;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B = CLBLM_L_X94Y126_SLICE_X149Y126_BO6;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C = CLBLM_L_X94Y126_SLICE_X149Y126_CO6;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D = CLBLM_L_X94Y126_SLICE_X149Y126_DO6;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A = CLBLM_L_X94Y127_SLICE_X148Y127_AO6;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B = CLBLM_L_X94Y127_SLICE_X148Y127_BO6;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C = CLBLM_L_X94Y127_SLICE_X148Y127_CO6;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D = CLBLM_L_X94Y127_SLICE_X148Y127_DO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A = CLBLM_L_X94Y127_SLICE_X149Y127_AO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B = CLBLM_L_X94Y127_SLICE_X149Y127_BO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C = CLBLM_L_X94Y127_SLICE_X149Y127_CO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D = CLBLM_L_X94Y127_SLICE_X149Y127_DO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_AMUX = CLBLM_L_X94Y127_SLICE_X149Y127_A5Q;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_BMUX = CLBLM_L_X94Y127_SLICE_X149Y127_B5Q;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_CMUX = CLBLM_L_X94Y127_SLICE_X149Y127_CO5;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A = CLBLM_L_X94Y128_SLICE_X148Y128_AO6;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B = CLBLM_L_X94Y128_SLICE_X148Y128_BO6;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C = CLBLM_L_X94Y128_SLICE_X148Y128_CO6;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D = CLBLM_L_X94Y128_SLICE_X148Y128_DO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A = CLBLM_L_X94Y128_SLICE_X149Y128_AO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B = CLBLM_L_X94Y128_SLICE_X149Y128_BO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C = CLBLM_L_X94Y128_SLICE_X149Y128_CO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D = CLBLM_L_X94Y128_SLICE_X149Y128_DO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_AMUX = CLBLM_L_X94Y128_SLICE_X149Y128_A5Q;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_BMUX = CLBLM_L_X94Y128_SLICE_X149Y128_BO5;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_CMUX = CLBLM_L_X94Y128_SLICE_X149Y128_C5Q;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A = CLBLM_L_X94Y129_SLICE_X148Y129_AO6;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B = CLBLM_L_X94Y129_SLICE_X148Y129_BO6;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C = CLBLM_L_X94Y129_SLICE_X148Y129_CO6;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D = CLBLM_L_X94Y129_SLICE_X148Y129_DO6;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_BMUX = CLBLM_L_X94Y129_SLICE_X148Y129_B5Q;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A = CLBLM_L_X94Y129_SLICE_X149Y129_AO6;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B = CLBLM_L_X94Y129_SLICE_X149Y129_BO6;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C = CLBLM_L_X94Y129_SLICE_X149Y129_CO6;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D = CLBLM_L_X94Y129_SLICE_X149Y129_DO6;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A = CLBLM_L_X94Y130_SLICE_X148Y130_AO6;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B = CLBLM_L_X94Y130_SLICE_X148Y130_BO6;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C = CLBLM_L_X94Y130_SLICE_X148Y130_CO6;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D = CLBLM_L_X94Y130_SLICE_X148Y130_DO6;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A = CLBLM_L_X94Y130_SLICE_X149Y130_AO6;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B = CLBLM_L_X94Y130_SLICE_X149Y130_BO6;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C = CLBLM_L_X94Y130_SLICE_X149Y130_CO6;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D = CLBLM_L_X94Y130_SLICE_X149Y130_DO6;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_AMUX = CLBLM_L_X94Y130_SLICE_X149Y130_A5Q;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A = CLBLM_L_X94Y132_SLICE_X148Y132_AO6;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B = CLBLM_L_X94Y132_SLICE_X148Y132_BO6;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C = CLBLM_L_X94Y132_SLICE_X148Y132_CO6;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D = CLBLM_L_X94Y132_SLICE_X148Y132_DO6;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A = CLBLM_L_X94Y132_SLICE_X149Y132_AO6;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B = CLBLM_L_X94Y132_SLICE_X149Y132_BO6;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C = CLBLM_L_X94Y132_SLICE_X149Y132_CO6;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D = CLBLM_L_X94Y132_SLICE_X149Y132_DO6;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_AMUX = CLBLM_L_X94Y132_SLICE_X149Y132_AO6;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A = CLBLM_L_X98Y110_SLICE_X154Y110_AO6;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B = CLBLM_L_X98Y110_SLICE_X154Y110_BO6;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C = CLBLM_L_X98Y110_SLICE_X154Y110_CO6;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D = CLBLM_L_X98Y110_SLICE_X154Y110_DO6;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_AMUX = CLBLM_L_X98Y110_SLICE_X154Y110_A5Q;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A = CLBLM_L_X98Y110_SLICE_X155Y110_AO6;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B = CLBLM_L_X98Y110_SLICE_X155Y110_BO6;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C = CLBLM_L_X98Y110_SLICE_X155Y110_CO6;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D = CLBLM_L_X98Y110_SLICE_X155Y110_DO6;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A = CLBLM_L_X98Y111_SLICE_X154Y111_AO6;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B = CLBLM_L_X98Y111_SLICE_X154Y111_BO6;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C = CLBLM_L_X98Y111_SLICE_X154Y111_CO6;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D = CLBLM_L_X98Y111_SLICE_X154Y111_DO6;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_AMUX = CLBLM_L_X98Y111_SLICE_X154Y111_A5Q;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_BMUX = CLBLM_L_X98Y111_SLICE_X154Y111_B5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A = CLBLM_L_X98Y111_SLICE_X155Y111_AO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B = CLBLM_L_X98Y111_SLICE_X155Y111_BO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C = CLBLM_L_X98Y111_SLICE_X155Y111_CO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D = CLBLM_L_X98Y111_SLICE_X155Y111_DO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_AMUX = CLBLM_L_X98Y111_SLICE_X155Y111_A5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_BMUX = CLBLM_L_X98Y111_SLICE_X155Y111_B5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_CMUX = CLBLM_L_X98Y111_SLICE_X155Y111_C5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_DMUX = CLBLM_L_X98Y111_SLICE_X155Y111_DO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A = CLBLM_L_X98Y112_SLICE_X154Y112_AO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B = CLBLM_L_X98Y112_SLICE_X154Y112_BO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C = CLBLM_L_X98Y112_SLICE_X154Y112_CO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D = CLBLM_L_X98Y112_SLICE_X154Y112_DO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_AMUX = CLBLM_L_X98Y112_SLICE_X154Y112_A5Q;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_BMUX = CLBLM_L_X98Y112_SLICE_X154Y112_B5Q;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_CMUX = CLBLM_L_X98Y112_SLICE_X154Y112_CO6;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A = CLBLM_L_X98Y112_SLICE_X155Y112_AO6;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B = CLBLM_L_X98Y112_SLICE_X155Y112_BO6;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C = CLBLM_L_X98Y112_SLICE_X155Y112_CO6;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D = CLBLM_L_X98Y112_SLICE_X155Y112_DO6;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_AMUX = CLBLM_L_X98Y112_SLICE_X155Y112_A5Q;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A = CLBLM_L_X98Y113_SLICE_X154Y113_AO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B = CLBLM_L_X98Y113_SLICE_X154Y113_BO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C = CLBLM_L_X98Y113_SLICE_X154Y113_CO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D = CLBLM_L_X98Y113_SLICE_X154Y113_DO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_AMUX = CLBLM_L_X98Y113_SLICE_X154Y113_A5Q;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A = CLBLM_L_X98Y113_SLICE_X155Y113_AO6;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B = CLBLM_L_X98Y113_SLICE_X155Y113_BO6;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C = CLBLM_L_X98Y113_SLICE_X155Y113_CO6;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D = CLBLM_L_X98Y113_SLICE_X155Y113_DO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A = CLBLM_L_X98Y114_SLICE_X154Y114_AO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B = CLBLM_L_X98Y114_SLICE_X154Y114_BO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C = CLBLM_L_X98Y114_SLICE_X154Y114_CO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D = CLBLM_L_X98Y114_SLICE_X154Y114_DO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_AMUX = CLBLM_L_X98Y114_SLICE_X154Y114_A5Q;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_BMUX = CLBLM_L_X98Y114_SLICE_X154Y114_B5Q;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_CMUX = CLBLM_L_X98Y114_SLICE_X154Y114_C5Q;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A = CLBLM_L_X98Y114_SLICE_X155Y114_AO6;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B = CLBLM_L_X98Y114_SLICE_X155Y114_BO6;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C = CLBLM_L_X98Y114_SLICE_X155Y114_CO6;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D = CLBLM_L_X98Y114_SLICE_X155Y114_DO6;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A = CLBLM_L_X98Y115_SLICE_X154Y115_AO6;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B = CLBLM_L_X98Y115_SLICE_X154Y115_BO6;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C = CLBLM_L_X98Y115_SLICE_X154Y115_CO6;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D = CLBLM_L_X98Y115_SLICE_X154Y115_DO6;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_AMUX = CLBLM_L_X98Y115_SLICE_X154Y115_A5Q;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_BMUX = CLBLM_L_X98Y115_SLICE_X154Y115_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A = CLBLM_L_X98Y115_SLICE_X155Y115_AO6;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B = CLBLM_L_X98Y115_SLICE_X155Y115_BO6;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C = CLBLM_L_X98Y115_SLICE_X155Y115_CO6;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D = CLBLM_L_X98Y115_SLICE_X155Y115_DO6;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_AMUX = CLBLM_L_X98Y115_SLICE_X155Y115_A5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_BMUX = CLBLM_L_X98Y115_SLICE_X155Y115_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_CMUX = CLBLM_L_X98Y115_SLICE_X155Y115_C5Q;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A = CLBLM_L_X98Y116_SLICE_X154Y116_AO6;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B = CLBLM_L_X98Y116_SLICE_X154Y116_BO6;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C = CLBLM_L_X98Y116_SLICE_X154Y116_CO6;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D = CLBLM_L_X98Y116_SLICE_X154Y116_DO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A = CLBLM_L_X98Y116_SLICE_X155Y116_AO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B = CLBLM_L_X98Y116_SLICE_X155Y116_BO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C = CLBLM_L_X98Y116_SLICE_X155Y116_CO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D = CLBLM_L_X98Y116_SLICE_X155Y116_DO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_AMUX = CLBLM_L_X98Y116_SLICE_X155Y116_A5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_BMUX = CLBLM_L_X98Y116_SLICE_X155Y116_B5Q;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A = CLBLM_L_X98Y117_SLICE_X154Y117_AO6;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B = CLBLM_L_X98Y117_SLICE_X154Y117_BO6;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C = CLBLM_L_X98Y117_SLICE_X154Y117_CO6;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D = CLBLM_L_X98Y117_SLICE_X154Y117_DO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A = CLBLM_L_X98Y117_SLICE_X155Y117_AO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B = CLBLM_L_X98Y117_SLICE_X155Y117_BO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C = CLBLM_L_X98Y117_SLICE_X155Y117_CO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D = CLBLM_L_X98Y117_SLICE_X155Y117_DO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_AMUX = CLBLM_L_X98Y117_SLICE_X155Y117_A5Q;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_BMUX = CLBLM_L_X98Y117_SLICE_X155Y117_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A = CLBLM_L_X98Y119_SLICE_X154Y119_AO6;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B = CLBLM_L_X98Y119_SLICE_X154Y119_BO6;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C = CLBLM_L_X98Y119_SLICE_X154Y119_CO6;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D = CLBLM_L_X98Y119_SLICE_X154Y119_DO6;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_AMUX = CLBLM_L_X98Y119_SLICE_X154Y119_A5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_BMUX = CLBLM_L_X98Y119_SLICE_X154Y119_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_CMUX = CLBLM_L_X98Y119_SLICE_X154Y119_CO5;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A = CLBLM_L_X98Y119_SLICE_X155Y119_AO6;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B = CLBLM_L_X98Y119_SLICE_X155Y119_BO6;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C = CLBLM_L_X98Y119_SLICE_X155Y119_CO6;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D = CLBLM_L_X98Y119_SLICE_X155Y119_DO6;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_BMUX = CLBLM_L_X98Y119_SLICE_X155Y119_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_CMUX = CLBLM_L_X98Y119_SLICE_X155Y119_C5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A = CLBLM_L_X98Y120_SLICE_X154Y120_AO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B = CLBLM_L_X98Y120_SLICE_X154Y120_BO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C = CLBLM_L_X98Y120_SLICE_X154Y120_CO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D = CLBLM_L_X98Y120_SLICE_X154Y120_DO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_AMUX = CLBLM_L_X98Y120_SLICE_X154Y120_A5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_BMUX = CLBLM_L_X98Y120_SLICE_X154Y120_BO5;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_CMUX = CLBLM_L_X98Y120_SLICE_X154Y120_C5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_DMUX = CLBLM_L_X98Y120_SLICE_X154Y120_DO6;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A = CLBLM_L_X98Y120_SLICE_X155Y120_AO6;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B = CLBLM_L_X98Y120_SLICE_X155Y120_BO6;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C = CLBLM_L_X98Y120_SLICE_X155Y120_CO6;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D = CLBLM_L_X98Y120_SLICE_X155Y120_DO6;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_AMUX = CLBLM_L_X98Y120_SLICE_X155Y120_A5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_BMUX = CLBLM_L_X98Y120_SLICE_X155Y120_B5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_DMUX = CLBLM_L_X98Y120_SLICE_X155Y120_DO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A = CLBLM_L_X98Y121_SLICE_X154Y121_AO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B = CLBLM_L_X98Y121_SLICE_X154Y121_BO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C = CLBLM_L_X98Y121_SLICE_X154Y121_CO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D = CLBLM_L_X98Y121_SLICE_X154Y121_DO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_AMUX = CLBLM_L_X98Y121_SLICE_X154Y121_A5Q;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_DMUX = CLBLM_L_X98Y121_SLICE_X154Y121_D5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A = CLBLM_L_X98Y121_SLICE_X155Y121_AO6;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B = CLBLM_L_X98Y121_SLICE_X155Y121_BO6;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C = CLBLM_L_X98Y121_SLICE_X155Y121_CO6;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D = CLBLM_L_X98Y121_SLICE_X155Y121_DO6;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_BMUX = CLBLM_L_X98Y121_SLICE_X155Y121_B5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_CMUX = CLBLM_L_X98Y121_SLICE_X155Y121_C5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A = CLBLM_L_X98Y122_SLICE_X154Y122_AO6;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B = CLBLM_L_X98Y122_SLICE_X154Y122_BO6;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C = CLBLM_L_X98Y122_SLICE_X154Y122_CO6;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D = CLBLM_L_X98Y122_SLICE_X154Y122_DO6;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_AMUX = CLBLM_L_X98Y122_SLICE_X154Y122_A5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_BMUX = CLBLM_L_X98Y122_SLICE_X154Y122_B5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A = CLBLM_L_X98Y122_SLICE_X155Y122_AO6;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B = CLBLM_L_X98Y122_SLICE_X155Y122_BO6;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C = CLBLM_L_X98Y122_SLICE_X155Y122_CO6;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D = CLBLM_L_X98Y122_SLICE_X155Y122_DO6;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_AMUX = CLBLM_L_X98Y122_SLICE_X155Y122_A5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_BMUX = CLBLM_L_X98Y122_SLICE_X155Y122_B5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A = CLBLM_L_X98Y123_SLICE_X154Y123_AO6;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B = CLBLM_L_X98Y123_SLICE_X154Y123_BO6;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C = CLBLM_L_X98Y123_SLICE_X154Y123_CO6;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D = CLBLM_L_X98Y123_SLICE_X154Y123_DO6;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_AMUX = CLBLM_L_X98Y123_SLICE_X154Y123_A5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_BMUX = CLBLM_L_X98Y123_SLICE_X154Y123_BO5;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_CMUX = CLBLM_L_X98Y123_SLICE_X154Y123_C5Q;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A = CLBLM_L_X98Y123_SLICE_X155Y123_AO6;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B = CLBLM_L_X98Y123_SLICE_X155Y123_BO6;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C = CLBLM_L_X98Y123_SLICE_X155Y123_CO6;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D = CLBLM_L_X98Y123_SLICE_X155Y123_DO6;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_AMUX = CLBLM_L_X98Y123_SLICE_X155Y123_A5Q;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_BMUX = CLBLM_L_X98Y123_SLICE_X155Y123_BO5;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_CMUX = CLBLM_L_X98Y123_SLICE_X155Y123_C5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A = CLBLM_L_X98Y124_SLICE_X154Y124_AO6;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B = CLBLM_L_X98Y124_SLICE_X154Y124_BO6;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C = CLBLM_L_X98Y124_SLICE_X154Y124_CO6;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D = CLBLM_L_X98Y124_SLICE_X154Y124_DO6;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_AMUX = CLBLM_L_X98Y124_SLICE_X154Y124_A5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_BMUX = CLBLM_L_X98Y124_SLICE_X154Y124_B5Q;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A = CLBLM_L_X98Y124_SLICE_X155Y124_AO6;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B = CLBLM_L_X98Y124_SLICE_X155Y124_BO6;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C = CLBLM_L_X98Y124_SLICE_X155Y124_CO6;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D = CLBLM_L_X98Y124_SLICE_X155Y124_DO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A = CLBLM_L_X98Y125_SLICE_X154Y125_AO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B = CLBLM_L_X98Y125_SLICE_X154Y125_BO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C = CLBLM_L_X98Y125_SLICE_X154Y125_CO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D = CLBLM_L_X98Y125_SLICE_X154Y125_DO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_AMUX = CLBLM_L_X98Y125_SLICE_X154Y125_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_BMUX = CLBLM_L_X98Y125_SLICE_X154Y125_B5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_CMUX = CLBLM_L_X98Y125_SLICE_X154Y125_C5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_DMUX = CLBLM_L_X98Y125_SLICE_X154Y125_D5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A = CLBLM_L_X98Y125_SLICE_X155Y125_AO6;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B = CLBLM_L_X98Y125_SLICE_X155Y125_BO6;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C = CLBLM_L_X98Y125_SLICE_X155Y125_CO6;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D = CLBLM_L_X98Y125_SLICE_X155Y125_DO6;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_AMUX = CLBLM_L_X98Y125_SLICE_X155Y125_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_BMUX = CLBLM_L_X98Y125_SLICE_X155Y125_BO5;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_CMUX = CLBLM_L_X98Y125_SLICE_X155Y125_C5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_DMUX = CLBLM_L_X98Y125_SLICE_X155Y125_DO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A = CLBLM_L_X98Y126_SLICE_X154Y126_AO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B = CLBLM_L_X98Y126_SLICE_X154Y126_BO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C = CLBLM_L_X98Y126_SLICE_X154Y126_CO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D = CLBLM_L_X98Y126_SLICE_X154Y126_DO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_AMUX = CLBLM_L_X98Y126_SLICE_X154Y126_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_BMUX = CLBLM_L_X98Y126_SLICE_X154Y126_B5Q;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_CMUX = CLBLM_L_X98Y126_SLICE_X154Y126_CO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A = CLBLM_L_X98Y126_SLICE_X155Y126_AO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B = CLBLM_L_X98Y126_SLICE_X155Y126_BO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C = CLBLM_L_X98Y126_SLICE_X155Y126_CO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D = CLBLM_L_X98Y126_SLICE_X155Y126_DO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_AMUX = CLBLM_L_X98Y126_SLICE_X155Y126_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_BMUX = CLBLM_L_X98Y126_SLICE_X155Y126_BO5;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_CMUX = CLBLM_L_X98Y126_SLICE_X155Y126_C5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A = CLBLM_L_X98Y127_SLICE_X154Y127_AO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B = CLBLM_L_X98Y127_SLICE_X154Y127_BO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C = CLBLM_L_X98Y127_SLICE_X154Y127_CO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D = CLBLM_L_X98Y127_SLICE_X154Y127_DO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_AMUX = CLBLM_L_X98Y127_SLICE_X154Y127_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_BMUX = CLBLM_L_X98Y127_SLICE_X154Y127_B5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_CMUX = CLBLM_L_X98Y127_SLICE_X154Y127_CO6;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A = CLBLM_L_X98Y127_SLICE_X155Y127_AO6;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B = CLBLM_L_X98Y127_SLICE_X155Y127_BO6;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C = CLBLM_L_X98Y127_SLICE_X155Y127_CO6;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D = CLBLM_L_X98Y127_SLICE_X155Y127_DO6;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_AMUX = CLBLM_L_X98Y127_SLICE_X155Y127_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_BMUX = CLBLM_L_X98Y127_SLICE_X155Y127_B5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A = CLBLM_L_X98Y128_SLICE_X154Y128_AO6;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B = CLBLM_L_X98Y128_SLICE_X154Y128_BO6;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C = CLBLM_L_X98Y128_SLICE_X154Y128_CO6;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D = CLBLM_L_X98Y128_SLICE_X154Y128_DO6;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_AMUX = CLBLM_L_X98Y128_SLICE_X154Y128_A5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_BMUX = CLBLM_L_X98Y128_SLICE_X154Y128_B5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_CMUX = CLBLM_L_X98Y128_SLICE_X154Y128_C5Q;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A = CLBLM_L_X98Y128_SLICE_X155Y128_AO6;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B = CLBLM_L_X98Y128_SLICE_X155Y128_BO6;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C = CLBLM_L_X98Y128_SLICE_X155Y128_CO6;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D = CLBLM_L_X98Y128_SLICE_X155Y128_DO6;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A = CLBLM_L_X98Y129_SLICE_X154Y129_AO6;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B = CLBLM_L_X98Y129_SLICE_X154Y129_BO6;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C = CLBLM_L_X98Y129_SLICE_X154Y129_CO6;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D = CLBLM_L_X98Y129_SLICE_X154Y129_DO6;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_AMUX = CLBLM_L_X98Y129_SLICE_X154Y129_AO5;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_BMUX = CLBLM_L_X98Y129_SLICE_X154Y129_B5Q;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A = CLBLM_L_X98Y129_SLICE_X155Y129_AO6;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B = CLBLM_L_X98Y129_SLICE_X155Y129_BO6;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C = CLBLM_L_X98Y129_SLICE_X155Y129_CO6;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D = CLBLM_L_X98Y129_SLICE_X155Y129_DO6;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_AMUX = CLBLM_L_X98Y129_SLICE_X155Y129_A5Q;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_BMUX = CLBLM_L_X98Y129_SLICE_X155Y129_BO5;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_CMUX = CLBLM_L_X98Y129_SLICE_X155Y129_C5Q;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A = CLBLM_L_X98Y130_SLICE_X154Y130_AO6;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B = CLBLM_L_X98Y130_SLICE_X154Y130_BO6;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C = CLBLM_L_X98Y130_SLICE_X154Y130_CO6;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D = CLBLM_L_X98Y130_SLICE_X154Y130_DO6;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_AMUX = CLBLM_L_X98Y130_SLICE_X154Y130_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_BMUX = CLBLM_L_X98Y130_SLICE_X154Y130_BO5;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_CMUX = CLBLM_L_X98Y130_SLICE_X154Y130_C5Q;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A = CLBLM_L_X98Y130_SLICE_X155Y130_AO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B = CLBLM_L_X98Y130_SLICE_X155Y130_BO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C = CLBLM_L_X98Y130_SLICE_X155Y130_CO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D = CLBLM_L_X98Y130_SLICE_X155Y130_DO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_AMUX = CLBLM_L_X98Y130_SLICE_X155Y130_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_DMUX = CLBLM_L_X98Y130_SLICE_X155Y130_D5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B = CLBLM_L_X98Y131_SLICE_X154Y131_BO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C = CLBLM_L_X98Y131_SLICE_X154Y131_CO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D = CLBLM_L_X98Y131_SLICE_X154Y131_DO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_AMUX = CLBLM_L_X98Y131_SLICE_X154Y131_A5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_BMUX = CLBLM_L_X98Y131_SLICE_X154Y131_BO5;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_CMUX = CLBLM_L_X98Y131_SLICE_X154Y131_C5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A = CLBLM_L_X98Y131_SLICE_X155Y131_AO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B = CLBLM_L_X98Y131_SLICE_X155Y131_BO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C = CLBLM_L_X98Y131_SLICE_X155Y131_CO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D = CLBLM_L_X98Y131_SLICE_X155Y131_DO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_AMUX = CLBLM_L_X98Y131_SLICE_X155Y131_A5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_BMUX = CLBLM_L_X98Y131_SLICE_X155Y131_B5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_CMUX = CLBLM_L_X98Y131_SLICE_X155Y131_CO5;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_DMUX = CLBLM_L_X98Y131_SLICE_X155Y131_D5Q;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B = CLBLM_L_X98Y132_SLICE_X154Y132_BO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C = CLBLM_L_X98Y132_SLICE_X154Y132_CO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D = CLBLM_L_X98Y132_SLICE_X154Y132_DO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_AMUX = CLBLM_L_X98Y132_SLICE_X154Y132_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_BMUX = CLBLM_L_X98Y132_SLICE_X154Y132_BO5;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_CMUX = CLBLM_L_X98Y132_SLICE_X154Y132_C5Q;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A = CLBLM_L_X98Y132_SLICE_X155Y132_AO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B = CLBLM_L_X98Y132_SLICE_X155Y132_BO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C = CLBLM_L_X98Y132_SLICE_X155Y132_CO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D = CLBLM_L_X98Y132_SLICE_X155Y132_DO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_CMUX = CLBLM_L_X98Y132_SLICE_X155Y132_C5Q;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A = CLBLM_L_X98Y133_SLICE_X154Y133_AO6;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B = CLBLM_L_X98Y133_SLICE_X154Y133_BO6;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C = CLBLM_L_X98Y133_SLICE_X154Y133_CO6;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D = CLBLM_L_X98Y133_SLICE_X154Y133_DO6;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_AMUX = CLBLM_L_X98Y133_SLICE_X154Y133_A5Q;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_BMUX = CLBLM_L_X98Y133_SLICE_X154Y133_B5Q;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A = CLBLM_L_X98Y133_SLICE_X155Y133_AO6;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B = CLBLM_L_X98Y133_SLICE_X155Y133_BO6;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C = CLBLM_L_X98Y133_SLICE_X155Y133_CO6;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D = CLBLM_L_X98Y133_SLICE_X155Y133_DO6;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_AMUX = CLBLM_L_X98Y133_SLICE_X155Y133_A5Q;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A = CLBLM_L_X98Y134_SLICE_X154Y134_AO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B = CLBLM_L_X98Y134_SLICE_X154Y134_BO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C = CLBLM_L_X98Y134_SLICE_X154Y134_CO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D = CLBLM_L_X98Y134_SLICE_X154Y134_DO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_AMUX = CLBLM_L_X98Y134_SLICE_X154Y134_A5Q;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_BMUX = CLBLM_L_X98Y134_SLICE_X154Y134_BO5;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_CMUX = CLBLM_L_X98Y134_SLICE_X154Y134_C5Q;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A = CLBLM_L_X98Y134_SLICE_X155Y134_AO6;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B = CLBLM_L_X98Y134_SLICE_X155Y134_BO6;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C = CLBLM_L_X98Y134_SLICE_X155Y134_CO6;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D = CLBLM_L_X98Y134_SLICE_X155Y134_DO6;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A = CLBLM_R_X89Y114_SLICE_X140Y114_AO6;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B = CLBLM_R_X89Y114_SLICE_X140Y114_BO6;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C = CLBLM_R_X89Y114_SLICE_X140Y114_CO6;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D = CLBLM_R_X89Y114_SLICE_X140Y114_DO6;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A = CLBLM_R_X89Y114_SLICE_X141Y114_AO6;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B = CLBLM_R_X89Y114_SLICE_X141Y114_BO6;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C = CLBLM_R_X89Y114_SLICE_X141Y114_CO6;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D = CLBLM_R_X89Y114_SLICE_X141Y114_DO6;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_AMUX = CLBLM_R_X89Y114_SLICE_X141Y114_A5Q;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_BMUX = CLBLM_R_X89Y114_SLICE_X141Y114_B5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A = CLBLM_R_X89Y115_SLICE_X140Y115_AO6;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B = CLBLM_R_X89Y115_SLICE_X140Y115_BO6;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C = CLBLM_R_X89Y115_SLICE_X140Y115_CO6;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D = CLBLM_R_X89Y115_SLICE_X140Y115_DO6;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_AMUX = CLBLM_R_X89Y115_SLICE_X140Y115_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_BMUX = CLBLM_R_X89Y115_SLICE_X140Y115_BO5;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_CMUX = CLBLM_R_X89Y115_SLICE_X140Y115_C5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A = CLBLM_R_X89Y115_SLICE_X141Y115_AO6;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B = CLBLM_R_X89Y115_SLICE_X141Y115_BO6;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C = CLBLM_R_X89Y115_SLICE_X141Y115_CO6;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D = CLBLM_R_X89Y115_SLICE_X141Y115_DO6;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_AMUX = CLBLM_R_X89Y115_SLICE_X141Y115_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_BMUX = CLBLM_R_X89Y115_SLICE_X141Y115_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A = CLBLM_R_X89Y116_SLICE_X140Y116_AO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B = CLBLM_R_X89Y116_SLICE_X140Y116_BO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C = CLBLM_R_X89Y116_SLICE_X140Y116_CO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D = CLBLM_R_X89Y116_SLICE_X140Y116_DO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_AMUX = CLBLM_R_X89Y116_SLICE_X140Y116_A5Q;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_BMUX = CLBLM_R_X89Y116_SLICE_X140Y116_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A = CLBLM_R_X89Y116_SLICE_X141Y116_AO6;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B = CLBLM_R_X89Y116_SLICE_X141Y116_BO6;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C = CLBLM_R_X89Y116_SLICE_X141Y116_CO6;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D = CLBLM_R_X89Y116_SLICE_X141Y116_DO6;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_AMUX = CLBLM_R_X89Y116_SLICE_X141Y116_AO5;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_BMUX = CLBLM_R_X89Y116_SLICE_X141Y116_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_CMUX = CLBLM_R_X89Y116_SLICE_X141Y116_C5Q;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A = CLBLM_R_X89Y117_SLICE_X140Y117_AO6;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B = CLBLM_R_X89Y117_SLICE_X140Y117_BO6;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C = CLBLM_R_X89Y117_SLICE_X140Y117_CO6;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D = CLBLM_R_X89Y117_SLICE_X140Y117_DO6;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_AMUX = CLBLM_R_X89Y117_SLICE_X140Y117_A5Q;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_CMUX = CLBLM_R_X89Y117_SLICE_X140Y117_C5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A = CLBLM_R_X89Y117_SLICE_X141Y117_AO6;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B = CLBLM_R_X89Y117_SLICE_X141Y117_BO6;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C = CLBLM_R_X89Y117_SLICE_X141Y117_CO6;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D = CLBLM_R_X89Y117_SLICE_X141Y117_DO6;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_AMUX = CLBLM_R_X89Y117_SLICE_X141Y117_A5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_BMUX = CLBLM_R_X89Y117_SLICE_X141Y117_BO5;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_CMUX = CLBLM_R_X89Y117_SLICE_X141Y117_C5Q;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A = CLBLM_R_X89Y118_SLICE_X140Y118_AO6;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B = CLBLM_R_X89Y118_SLICE_X140Y118_BO6;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C = CLBLM_R_X89Y118_SLICE_X140Y118_CO6;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D = CLBLM_R_X89Y118_SLICE_X140Y118_DO6;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_AMUX = CLBLM_R_X89Y118_SLICE_X140Y118_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_BMUX = CLBLM_R_X89Y118_SLICE_X140Y118_B5Q;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_CMUX = CLBLM_R_X89Y118_SLICE_X140Y118_CO5;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_DMUX = CLBLM_R_X89Y118_SLICE_X140Y118_D5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A = CLBLM_R_X89Y118_SLICE_X141Y118_AO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B = CLBLM_R_X89Y118_SLICE_X141Y118_BO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C = CLBLM_R_X89Y118_SLICE_X141Y118_CO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D = CLBLM_R_X89Y118_SLICE_X141Y118_DO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_AMUX = CLBLM_R_X89Y118_SLICE_X141Y118_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_BMUX = CLBLM_R_X89Y118_SLICE_X141Y118_BO5;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_DMUX = CLBLM_R_X89Y118_SLICE_X141Y118_D5Q;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A = CLBLM_R_X89Y119_SLICE_X140Y119_AO6;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B = CLBLM_R_X89Y119_SLICE_X140Y119_BO6;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C = CLBLM_R_X89Y119_SLICE_X140Y119_CO6;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D = CLBLM_R_X89Y119_SLICE_X140Y119_DO6;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_AMUX = CLBLM_R_X89Y119_SLICE_X140Y119_A5Q;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_BMUX = CLBLM_R_X89Y119_SLICE_X140Y119_B5Q;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A = CLBLM_R_X89Y119_SLICE_X141Y119_AO6;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B = CLBLM_R_X89Y119_SLICE_X141Y119_BO6;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C = CLBLM_R_X89Y119_SLICE_X141Y119_CO6;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D = CLBLM_R_X89Y119_SLICE_X141Y119_DO6;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_AMUX = CLBLM_R_X89Y119_SLICE_X141Y119_A5Q;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_BMUX = CLBLM_R_X89Y119_SLICE_X141Y119_BO5;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_CMUX = CLBLM_R_X89Y119_SLICE_X141Y119_C5Q;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A = CLBLM_R_X89Y120_SLICE_X140Y120_AO6;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B = CLBLM_R_X89Y120_SLICE_X140Y120_BO6;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C = CLBLM_R_X89Y120_SLICE_X140Y120_CO6;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D = CLBLM_R_X89Y120_SLICE_X140Y120_DO6;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_AMUX = CLBLM_R_X89Y120_SLICE_X140Y120_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_BMUX = CLBLM_R_X89Y120_SLICE_X140Y120_BO5;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A = CLBLM_R_X89Y120_SLICE_X141Y120_AO6;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B = CLBLM_R_X89Y120_SLICE_X141Y120_BO6;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C = CLBLM_R_X89Y120_SLICE_X141Y120_CO6;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D = CLBLM_R_X89Y120_SLICE_X141Y120_DO6;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_AMUX = CLBLM_R_X89Y120_SLICE_X141Y120_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_CMUX = CLBLM_R_X89Y120_SLICE_X141Y120_C5Q;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A = CLBLM_R_X89Y121_SLICE_X140Y121_AO6;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B = CLBLM_R_X89Y121_SLICE_X140Y121_BO6;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C = CLBLM_R_X89Y121_SLICE_X140Y121_CO6;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D = CLBLM_R_X89Y121_SLICE_X140Y121_DO6;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_AMUX = CLBLM_R_X89Y121_SLICE_X140Y121_A5Q;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_BMUX = CLBLM_R_X89Y121_SLICE_X140Y121_BO5;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_CMUX = CLBLM_R_X89Y121_SLICE_X140Y121_C5Q;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A = CLBLM_R_X89Y121_SLICE_X141Y121_AO6;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B = CLBLM_R_X89Y121_SLICE_X141Y121_BO6;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C = CLBLM_R_X89Y121_SLICE_X141Y121_CO6;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D = CLBLM_R_X89Y121_SLICE_X141Y121_DO6;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_AMUX = CLBLM_R_X89Y121_SLICE_X141Y121_A5Q;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_BMUX = CLBLM_R_X89Y121_SLICE_X141Y121_BO5;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_CMUX = CLBLM_R_X89Y121_SLICE_X141Y121_C5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A = CLBLM_R_X89Y122_SLICE_X140Y122_AO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B = CLBLM_R_X89Y122_SLICE_X140Y122_BO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C = CLBLM_R_X89Y122_SLICE_X140Y122_CO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D = CLBLM_R_X89Y122_SLICE_X140Y122_DO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_AMUX = CLBLM_R_X89Y122_SLICE_X140Y122_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_BMUX = CLBLM_R_X89Y122_SLICE_X140Y122_BO5;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_CMUX = CLBLM_R_X89Y122_SLICE_X140Y122_C5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A = CLBLM_R_X89Y122_SLICE_X141Y122_AO6;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B = CLBLM_R_X89Y122_SLICE_X141Y122_BO6;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C = CLBLM_R_X89Y122_SLICE_X141Y122_CO6;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D = CLBLM_R_X89Y122_SLICE_X141Y122_DO6;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_AMUX = CLBLM_R_X89Y122_SLICE_X141Y122_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_BMUX = CLBLM_R_X89Y122_SLICE_X141Y122_B5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_CMUX = CLBLM_R_X89Y122_SLICE_X141Y122_CO5;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_DMUX = CLBLM_R_X89Y122_SLICE_X141Y122_D5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A = CLBLM_R_X89Y123_SLICE_X140Y123_AO6;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B = CLBLM_R_X89Y123_SLICE_X140Y123_BO6;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C = CLBLM_R_X89Y123_SLICE_X140Y123_CO6;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D = CLBLM_R_X89Y123_SLICE_X140Y123_DO6;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_AMUX = CLBLM_R_X89Y123_SLICE_X140Y123_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_BMUX = CLBLM_R_X89Y123_SLICE_X140Y123_BO5;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_CMUX = CLBLM_R_X89Y123_SLICE_X140Y123_C5Q;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A = CLBLM_R_X89Y123_SLICE_X141Y123_AO6;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B = CLBLM_R_X89Y123_SLICE_X141Y123_BO6;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C = CLBLM_R_X89Y123_SLICE_X141Y123_CO6;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D = CLBLM_R_X89Y123_SLICE_X141Y123_DO6;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_AMUX = CLBLM_R_X89Y123_SLICE_X141Y123_A5Q;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A = CLBLM_R_X89Y124_SLICE_X140Y124_AO6;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B = CLBLM_R_X89Y124_SLICE_X140Y124_BO6;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C = CLBLM_R_X89Y124_SLICE_X140Y124_CO6;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D = CLBLM_R_X89Y124_SLICE_X140Y124_DO6;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_AMUX = CLBLM_R_X89Y124_SLICE_X140Y124_A5Q;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A = CLBLM_R_X89Y124_SLICE_X141Y124_AO6;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B = CLBLM_R_X89Y124_SLICE_X141Y124_BO6;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C = CLBLM_R_X89Y124_SLICE_X141Y124_CO6;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D = CLBLM_R_X89Y124_SLICE_X141Y124_DO6;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_AMUX = CLBLM_R_X89Y124_SLICE_X141Y124_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A = CLBLM_R_X89Y125_SLICE_X140Y125_AO6;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B = CLBLM_R_X89Y125_SLICE_X140Y125_BO6;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C = CLBLM_R_X89Y125_SLICE_X140Y125_CO6;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D = CLBLM_R_X89Y125_SLICE_X140Y125_DO6;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_AMUX = CLBLM_R_X89Y125_SLICE_X140Y125_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_BMUX = CLBLM_R_X89Y125_SLICE_X140Y125_B5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_CMUX = CLBLM_R_X89Y125_SLICE_X140Y125_CO5;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_DMUX = CLBLM_R_X89Y125_SLICE_X140Y125_D5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A = CLBLM_R_X89Y125_SLICE_X141Y125_AO6;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B = CLBLM_R_X89Y125_SLICE_X141Y125_BO6;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C = CLBLM_R_X89Y125_SLICE_X141Y125_CO6;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D = CLBLM_R_X89Y125_SLICE_X141Y125_DO6;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_AMUX = CLBLM_R_X89Y125_SLICE_X141Y125_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_BMUX = CLBLM_R_X89Y125_SLICE_X141Y125_BO5;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_CMUX = CLBLM_R_X89Y125_SLICE_X141Y125_C5Q;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A = CLBLM_R_X89Y126_SLICE_X140Y126_AO6;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B = CLBLM_R_X89Y126_SLICE_X140Y126_BO6;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C = CLBLM_R_X89Y126_SLICE_X140Y126_CO6;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D = CLBLM_R_X89Y126_SLICE_X140Y126_DO6;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_BMUX = CLBLM_R_X89Y126_SLICE_X140Y126_B5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A = CLBLM_R_X89Y126_SLICE_X141Y126_AO6;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B = CLBLM_R_X89Y126_SLICE_X141Y126_BO6;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C = CLBLM_R_X89Y126_SLICE_X141Y126_CO6;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D = CLBLM_R_X89Y126_SLICE_X141Y126_DO6;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_AMUX = CLBLM_R_X89Y126_SLICE_X141Y126_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_BMUX = CLBLM_R_X89Y126_SLICE_X141Y126_BO5;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_CMUX = CLBLM_R_X89Y126_SLICE_X141Y126_C5Q;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A = CLBLM_R_X89Y127_SLICE_X140Y127_AO6;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B = CLBLM_R_X89Y127_SLICE_X140Y127_BO6;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C = CLBLM_R_X89Y127_SLICE_X140Y127_CO6;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D = CLBLM_R_X89Y127_SLICE_X140Y127_DO6;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A = CLBLM_R_X89Y127_SLICE_X141Y127_AO6;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B = CLBLM_R_X89Y127_SLICE_X141Y127_BO6;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C = CLBLM_R_X89Y127_SLICE_X141Y127_CO6;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D = CLBLM_R_X89Y127_SLICE_X141Y127_DO6;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_AMUX = CLBLM_R_X89Y127_SLICE_X141Y127_A5Q;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A = CLBLM_R_X89Y128_SLICE_X140Y128_AO6;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B = CLBLM_R_X89Y128_SLICE_X140Y128_BO6;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C = CLBLM_R_X89Y128_SLICE_X140Y128_CO6;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D = CLBLM_R_X89Y128_SLICE_X140Y128_DO6;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_AMUX = CLBLM_R_X89Y128_SLICE_X140Y128_A5Q;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_BMUX = CLBLM_R_X89Y128_SLICE_X140Y128_BO5;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_CMUX = CLBLM_R_X89Y128_SLICE_X140Y128_C5Q;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A = CLBLM_R_X89Y128_SLICE_X141Y128_AO6;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B = CLBLM_R_X89Y128_SLICE_X141Y128_BO6;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C = CLBLM_R_X89Y128_SLICE_X141Y128_CO6;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D = CLBLM_R_X89Y128_SLICE_X141Y128_DO6;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_AMUX = CLBLM_R_X89Y128_SLICE_X141Y128_A5Q;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A = CLBLM_R_X89Y130_SLICE_X140Y130_AO6;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B = CLBLM_R_X89Y130_SLICE_X140Y130_BO6;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C = CLBLM_R_X89Y130_SLICE_X140Y130_CO6;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D = CLBLM_R_X89Y130_SLICE_X140Y130_DO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A = CLBLM_R_X89Y130_SLICE_X141Y130_AO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B = CLBLM_R_X89Y130_SLICE_X141Y130_BO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C = CLBLM_R_X89Y130_SLICE_X141Y130_CO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D = CLBLM_R_X89Y130_SLICE_X141Y130_DO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_AMUX = CLBLM_R_X89Y130_SLICE_X141Y130_A5Q;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A = CLBLM_R_X89Y131_SLICE_X140Y131_AO6;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B = CLBLM_R_X89Y131_SLICE_X140Y131_BO6;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C = CLBLM_R_X89Y131_SLICE_X140Y131_CO6;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D = CLBLM_R_X89Y131_SLICE_X140Y131_DO6;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_AMUX = CLBLM_R_X89Y131_SLICE_X140Y131_A5Q;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A = CLBLM_R_X89Y131_SLICE_X141Y131_AO6;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B = CLBLM_R_X89Y131_SLICE_X141Y131_BO6;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C = CLBLM_R_X89Y131_SLICE_X141Y131_CO6;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D = CLBLM_R_X89Y131_SLICE_X141Y131_DO6;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A = CLBLM_R_X93Y111_SLICE_X146Y111_AO6;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B = CLBLM_R_X93Y111_SLICE_X146Y111_BO6;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C = CLBLM_R_X93Y111_SLICE_X146Y111_CO6;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D = CLBLM_R_X93Y111_SLICE_X146Y111_DO6;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A = CLBLM_R_X93Y111_SLICE_X147Y111_AO6;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B = CLBLM_R_X93Y111_SLICE_X147Y111_BO6;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C = CLBLM_R_X93Y111_SLICE_X147Y111_CO6;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D = CLBLM_R_X93Y111_SLICE_X147Y111_DO6;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_AMUX = CLBLM_R_X93Y111_SLICE_X147Y111_A5Q;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_BMUX = CLBLM_R_X93Y111_SLICE_X147Y111_B5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A = CLBLM_R_X93Y112_SLICE_X146Y112_AO6;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B = CLBLM_R_X93Y112_SLICE_X146Y112_BO6;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C = CLBLM_R_X93Y112_SLICE_X146Y112_CO6;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D = CLBLM_R_X93Y112_SLICE_X146Y112_DO6;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_AMUX = CLBLM_R_X93Y112_SLICE_X146Y112_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_BMUX = CLBLM_R_X93Y112_SLICE_X146Y112_B5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A = CLBLM_R_X93Y112_SLICE_X147Y112_AO6;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B = CLBLM_R_X93Y112_SLICE_X147Y112_BO6;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C = CLBLM_R_X93Y112_SLICE_X147Y112_CO6;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D = CLBLM_R_X93Y112_SLICE_X147Y112_DO6;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_AMUX = CLBLM_R_X93Y112_SLICE_X147Y112_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_BMUX = CLBLM_R_X93Y112_SLICE_X147Y112_B5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_CMUX = CLBLM_R_X93Y112_SLICE_X147Y112_C5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A = CLBLM_R_X93Y113_SLICE_X146Y113_AO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B = CLBLM_R_X93Y113_SLICE_X146Y113_BO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C = CLBLM_R_X93Y113_SLICE_X146Y113_CO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D = CLBLM_R_X93Y113_SLICE_X146Y113_DO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_AMUX = CLBLM_R_X93Y113_SLICE_X146Y113_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_BMUX = CLBLM_R_X93Y113_SLICE_X146Y113_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A = CLBLM_R_X93Y113_SLICE_X147Y113_AO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B = CLBLM_R_X93Y113_SLICE_X147Y113_BO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C = CLBLM_R_X93Y113_SLICE_X147Y113_CO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D = CLBLM_R_X93Y113_SLICE_X147Y113_DO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_AMUX = CLBLM_R_X93Y113_SLICE_X147Y113_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_BMUX = CLBLM_R_X93Y113_SLICE_X147Y113_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A = CLBLM_R_X93Y114_SLICE_X146Y114_AO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B = CLBLM_R_X93Y114_SLICE_X146Y114_BO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C = CLBLM_R_X93Y114_SLICE_X146Y114_CO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D = CLBLM_R_X93Y114_SLICE_X146Y114_DO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_AMUX = CLBLM_R_X93Y114_SLICE_X146Y114_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_BMUX = CLBLM_R_X93Y114_SLICE_X146Y114_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_DMUX = CLBLM_R_X93Y114_SLICE_X146Y114_DO6;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A = CLBLM_R_X93Y114_SLICE_X147Y114_AO6;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B = CLBLM_R_X93Y114_SLICE_X147Y114_BO6;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C = CLBLM_R_X93Y114_SLICE_X147Y114_CO6;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D = CLBLM_R_X93Y114_SLICE_X147Y114_DO6;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_AMUX = CLBLM_R_X93Y114_SLICE_X147Y114_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_BMUX = CLBLM_R_X93Y114_SLICE_X147Y114_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A = CLBLM_R_X93Y115_SLICE_X146Y115_AO6;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B = CLBLM_R_X93Y115_SLICE_X146Y115_BO6;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C = CLBLM_R_X93Y115_SLICE_X146Y115_CO6;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D = CLBLM_R_X93Y115_SLICE_X146Y115_DO6;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_AMUX = CLBLM_R_X93Y115_SLICE_X146Y115_A5Q;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_BMUX = CLBLM_R_X93Y115_SLICE_X146Y115_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A = CLBLM_R_X93Y115_SLICE_X147Y115_AO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B = CLBLM_R_X93Y115_SLICE_X147Y115_BO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C = CLBLM_R_X93Y115_SLICE_X147Y115_CO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D = CLBLM_R_X93Y115_SLICE_X147Y115_DO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_AMUX = CLBLM_R_X93Y115_SLICE_X147Y115_A5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_BMUX = CLBLM_R_X93Y115_SLICE_X147Y115_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_CMUX = CLBLM_R_X93Y115_SLICE_X147Y115_CO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A = CLBLM_R_X93Y116_SLICE_X146Y116_AO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B = CLBLM_R_X93Y116_SLICE_X146Y116_BO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C = CLBLM_R_X93Y116_SLICE_X146Y116_CO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D = CLBLM_R_X93Y116_SLICE_X146Y116_DO6;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_AMUX = CLBLM_R_X93Y116_SLICE_X146Y116_A5Q;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_BMUX = CLBLM_R_X93Y116_SLICE_X146Y116_B5Q;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A = CLBLM_R_X93Y116_SLICE_X147Y116_AO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B = CLBLM_R_X93Y116_SLICE_X147Y116_BO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C = CLBLM_R_X93Y116_SLICE_X147Y116_CO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D = CLBLM_R_X93Y116_SLICE_X147Y116_DO6;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_AMUX = CLBLM_R_X93Y116_SLICE_X147Y116_A5Q;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_BMUX = CLBLM_R_X93Y116_SLICE_X147Y116_B5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A = CLBLM_R_X93Y117_SLICE_X146Y117_AO6;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B = CLBLM_R_X93Y117_SLICE_X146Y117_BO6;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C = CLBLM_R_X93Y117_SLICE_X146Y117_CO6;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D = CLBLM_R_X93Y117_SLICE_X146Y117_DO6;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_AMUX = CLBLM_R_X93Y117_SLICE_X146Y117_A5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_BMUX = CLBLM_R_X93Y117_SLICE_X146Y117_B5Q;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A = CLBLM_R_X93Y117_SLICE_X147Y117_AO6;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B = CLBLM_R_X93Y117_SLICE_X147Y117_BO6;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C = CLBLM_R_X93Y117_SLICE_X147Y117_CO6;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D = CLBLM_R_X93Y117_SLICE_X147Y117_DO6;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A = CLBLM_R_X93Y118_SLICE_X146Y118_AO6;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B = CLBLM_R_X93Y118_SLICE_X146Y118_BO6;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C = CLBLM_R_X93Y118_SLICE_X146Y118_CO6;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D = CLBLM_R_X93Y118_SLICE_X146Y118_DO6;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A = CLBLM_R_X93Y118_SLICE_X147Y118_AO6;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B = CLBLM_R_X93Y118_SLICE_X147Y118_BO6;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C = CLBLM_R_X93Y118_SLICE_X147Y118_CO6;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D = CLBLM_R_X93Y118_SLICE_X147Y118_DO6;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_AMUX = CLBLM_R_X93Y118_SLICE_X147Y118_A5Q;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_BMUX = CLBLM_R_X93Y118_SLICE_X147Y118_B5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A = CLBLM_R_X93Y119_SLICE_X146Y119_AO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B = CLBLM_R_X93Y119_SLICE_X146Y119_BO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C = CLBLM_R_X93Y119_SLICE_X146Y119_CO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D = CLBLM_R_X93Y119_SLICE_X146Y119_DO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_AMUX = CLBLM_R_X93Y119_SLICE_X146Y119_A5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_BMUX = CLBLM_R_X93Y119_SLICE_X146Y119_B5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_CMUX = CLBLM_R_X93Y119_SLICE_X146Y119_C5Q;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A = CLBLM_R_X93Y119_SLICE_X147Y119_AO6;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B = CLBLM_R_X93Y119_SLICE_X147Y119_BO6;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C = CLBLM_R_X93Y119_SLICE_X147Y119_CO6;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D = CLBLM_R_X93Y119_SLICE_X147Y119_DO6;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_AMUX = CLBLM_R_X93Y119_SLICE_X147Y119_A5Q;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_BMUX = CLBLM_R_X93Y119_SLICE_X147Y119_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A = CLBLM_R_X93Y120_SLICE_X146Y120_AO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B = CLBLM_R_X93Y120_SLICE_X146Y120_BO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C = CLBLM_R_X93Y120_SLICE_X146Y120_CO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D = CLBLM_R_X93Y120_SLICE_X146Y120_DO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_AMUX = CLBLM_R_X93Y120_SLICE_X146Y120_A5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_BMUX = CLBLM_R_X93Y120_SLICE_X146Y120_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A = CLBLM_R_X93Y120_SLICE_X147Y120_AO6;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B = CLBLM_R_X93Y120_SLICE_X147Y120_BO6;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C = CLBLM_R_X93Y120_SLICE_X147Y120_CO6;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D = CLBLM_R_X93Y120_SLICE_X147Y120_DO6;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_AMUX = CLBLM_R_X93Y120_SLICE_X147Y120_A5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_BMUX = CLBLM_R_X93Y120_SLICE_X147Y120_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_CMUX = CLBLM_R_X93Y120_SLICE_X147Y120_C5Q;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A = CLBLM_R_X93Y121_SLICE_X146Y121_AO6;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B = CLBLM_R_X93Y121_SLICE_X146Y121_BO6;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C = CLBLM_R_X93Y121_SLICE_X146Y121_CO6;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D = CLBLM_R_X93Y121_SLICE_X146Y121_DO6;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_AMUX = CLBLM_R_X93Y121_SLICE_X146Y121_A5Q;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A = CLBLM_R_X93Y121_SLICE_X147Y121_AO6;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B = CLBLM_R_X93Y121_SLICE_X147Y121_BO6;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C = CLBLM_R_X93Y121_SLICE_X147Y121_CO6;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D = CLBLM_R_X93Y121_SLICE_X147Y121_DO6;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_AMUX = CLBLM_R_X93Y121_SLICE_X147Y121_AO6;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_BMUX = CLBLM_R_X93Y121_SLICE_X147Y121_B5Q;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_CMUX = CLBLM_R_X93Y121_SLICE_X147Y121_C5Q;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A = CLBLM_R_X93Y122_SLICE_X146Y122_AO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B = CLBLM_R_X93Y122_SLICE_X146Y122_BO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C = CLBLM_R_X93Y122_SLICE_X146Y122_CO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D = CLBLM_R_X93Y122_SLICE_X146Y122_DO6;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_AMUX = CLBLM_R_X93Y122_SLICE_X146Y122_A5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A = CLBLM_R_X93Y122_SLICE_X147Y122_AO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B = CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C = CLBLM_R_X93Y122_SLICE_X147Y122_CO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D = CLBLM_R_X93Y122_SLICE_X147Y122_DO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_AMUX = CLBLM_R_X93Y122_SLICE_X147Y122_A5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_BMUX = CLBLM_R_X93Y122_SLICE_X147Y122_BO5;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_CMUX = CLBLM_R_X93Y122_SLICE_X147Y122_C5Q;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A = CLBLM_R_X93Y123_SLICE_X146Y123_AO6;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B = CLBLM_R_X93Y123_SLICE_X146Y123_BO6;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C = CLBLM_R_X93Y123_SLICE_X146Y123_CO6;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D = CLBLM_R_X93Y123_SLICE_X146Y123_DO6;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_BMUX = CLBLM_R_X93Y123_SLICE_X146Y123_B5Q;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A = CLBLM_R_X93Y123_SLICE_X147Y123_AO6;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B = CLBLM_R_X93Y123_SLICE_X147Y123_BO6;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C = CLBLM_R_X93Y123_SLICE_X147Y123_CO6;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D = CLBLM_R_X93Y123_SLICE_X147Y123_DO6;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_AMUX = CLBLM_R_X93Y123_SLICE_X147Y123_AO5;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_BMUX = CLBLM_R_X93Y123_SLICE_X147Y123_B5Q;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_CMUX = CLBLM_R_X93Y123_SLICE_X147Y123_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A = CLBLM_R_X93Y124_SLICE_X146Y124_AO6;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B = CLBLM_R_X93Y124_SLICE_X146Y124_BO6;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C = CLBLM_R_X93Y124_SLICE_X146Y124_CO6;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D = CLBLM_R_X93Y124_SLICE_X146Y124_DO6;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_AMUX = CLBLM_R_X93Y124_SLICE_X146Y124_A5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_BMUX = CLBLM_R_X93Y124_SLICE_X146Y124_BO5;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_CMUX = CLBLM_R_X93Y124_SLICE_X146Y124_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A = CLBLM_R_X93Y124_SLICE_X147Y124_AO6;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B = CLBLM_R_X93Y124_SLICE_X147Y124_BO6;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C = CLBLM_R_X93Y124_SLICE_X147Y124_CO6;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D = CLBLM_R_X93Y124_SLICE_X147Y124_DO6;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_AMUX = CLBLM_R_X93Y124_SLICE_X147Y124_A5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_BMUX = CLBLM_R_X93Y124_SLICE_X147Y124_B5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_CMUX = CLBLM_R_X93Y124_SLICE_X147Y124_C5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A = CLBLM_R_X93Y125_SLICE_X146Y125_AO6;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B = CLBLM_R_X93Y125_SLICE_X146Y125_BO6;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C = CLBLM_R_X93Y125_SLICE_X146Y125_CO6;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D = CLBLM_R_X93Y125_SLICE_X146Y125_DO6;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_AMUX = CLBLM_R_X93Y125_SLICE_X146Y125_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_BMUX = CLBLM_R_X93Y125_SLICE_X146Y125_BO5;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_CMUX = CLBLM_R_X93Y125_SLICE_X146Y125_C5Q;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A = CLBLM_R_X93Y125_SLICE_X147Y125_AO6;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B = CLBLM_R_X93Y125_SLICE_X147Y125_BO6;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C = CLBLM_R_X93Y125_SLICE_X147Y125_CO6;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D = CLBLM_R_X93Y125_SLICE_X147Y125_DO6;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_AMUX = CLBLM_R_X93Y125_SLICE_X147Y125_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A = CLBLM_R_X93Y126_SLICE_X146Y126_AO6;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B = CLBLM_R_X93Y126_SLICE_X146Y126_BO6;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C = CLBLM_R_X93Y126_SLICE_X146Y126_CO6;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D = CLBLM_R_X93Y126_SLICE_X146Y126_DO6;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_AMUX = CLBLM_R_X93Y126_SLICE_X146Y126_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_CMUX = CLBLM_R_X93Y126_SLICE_X146Y126_C5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A = CLBLM_R_X93Y126_SLICE_X147Y126_AO6;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B = CLBLM_R_X93Y126_SLICE_X147Y126_BO6;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C = CLBLM_R_X93Y126_SLICE_X147Y126_CO6;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D = CLBLM_R_X93Y126_SLICE_X147Y126_DO6;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_AMUX = CLBLM_R_X93Y126_SLICE_X147Y126_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_BMUX = CLBLM_R_X93Y126_SLICE_X147Y126_BO5;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_CMUX = CLBLM_R_X93Y126_SLICE_X147Y126_C5Q;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A = CLBLM_R_X93Y127_SLICE_X146Y127_AO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B = CLBLM_R_X93Y127_SLICE_X146Y127_BO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C = CLBLM_R_X93Y127_SLICE_X146Y127_CO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D = CLBLM_R_X93Y127_SLICE_X146Y127_DO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_AMUX = CLBLM_R_X93Y127_SLICE_X146Y127_A5Q;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A = CLBLM_R_X93Y127_SLICE_X147Y127_AO6;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B = CLBLM_R_X93Y127_SLICE_X147Y127_BO6;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C = CLBLM_R_X93Y127_SLICE_X147Y127_CO6;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D = CLBLM_R_X93Y127_SLICE_X147Y127_DO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A = CLBLM_R_X93Y128_SLICE_X146Y128_AO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B = CLBLM_R_X93Y128_SLICE_X146Y128_BO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C = CLBLM_R_X93Y128_SLICE_X146Y128_CO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D = CLBLM_R_X93Y128_SLICE_X146Y128_DO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_AMUX = CLBLM_R_X93Y128_SLICE_X146Y128_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_BMUX = CLBLM_R_X93Y128_SLICE_X146Y128_BO5;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_CMUX = CLBLM_R_X93Y128_SLICE_X146Y128_C5Q;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A = CLBLM_R_X93Y128_SLICE_X147Y128_AO6;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B = CLBLM_R_X93Y128_SLICE_X147Y128_BO6;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C = CLBLM_R_X93Y128_SLICE_X147Y128_CO6;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D = CLBLM_R_X93Y128_SLICE_X147Y128_DO6;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_AMUX = CLBLM_R_X93Y128_SLICE_X147Y128_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_BMUX = CLBLM_R_X93Y128_SLICE_X147Y128_B5Q;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A = CLBLM_R_X93Y129_SLICE_X146Y129_AO6;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B = CLBLM_R_X93Y129_SLICE_X146Y129_BO6;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C = CLBLM_R_X93Y129_SLICE_X146Y129_CO6;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D = CLBLM_R_X93Y129_SLICE_X146Y129_DO6;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_AMUX = CLBLM_R_X93Y129_SLICE_X146Y129_A5Q;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_BMUX = CLBLM_R_X93Y129_SLICE_X146Y129_B5Q;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A = CLBLM_R_X93Y129_SLICE_X147Y129_AO6;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B = CLBLM_R_X93Y129_SLICE_X147Y129_BO6;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C = CLBLM_R_X93Y129_SLICE_X147Y129_CO6;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D = CLBLM_R_X93Y129_SLICE_X147Y129_DO6;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_AMUX = CLBLM_R_X93Y129_SLICE_X147Y129_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A = CLBLM_R_X93Y130_SLICE_X146Y130_AO6;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B = CLBLM_R_X93Y130_SLICE_X146Y130_BO6;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C = CLBLM_R_X93Y130_SLICE_X146Y130_CO6;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D = CLBLM_R_X93Y130_SLICE_X146Y130_DO6;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_AMUX = CLBLM_R_X93Y130_SLICE_X146Y130_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_BMUX = CLBLM_R_X93Y130_SLICE_X146Y130_B5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A = CLBLM_R_X93Y130_SLICE_X147Y130_AO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B = CLBLM_R_X93Y130_SLICE_X147Y130_BO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C = CLBLM_R_X93Y130_SLICE_X147Y130_CO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D = CLBLM_R_X93Y130_SLICE_X147Y130_DO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_AMUX = CLBLM_R_X93Y130_SLICE_X147Y130_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_BMUX = CLBLM_R_X93Y130_SLICE_X147Y130_BO5;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_CMUX = CLBLM_R_X93Y130_SLICE_X147Y130_C5Q;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A = CLBLM_R_X93Y131_SLICE_X146Y131_AO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B = CLBLM_R_X93Y131_SLICE_X146Y131_BO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C = CLBLM_R_X93Y131_SLICE_X146Y131_CO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D = CLBLM_R_X93Y131_SLICE_X146Y131_DO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_AMUX = CLBLM_R_X93Y131_SLICE_X146Y131_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_BMUX = CLBLM_R_X93Y131_SLICE_X146Y131_BO5;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_CMUX = CLBLM_R_X93Y131_SLICE_X146Y131_C5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A = CLBLM_R_X93Y131_SLICE_X147Y131_AO6;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B = CLBLM_R_X93Y131_SLICE_X147Y131_BO6;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C = CLBLM_R_X93Y131_SLICE_X147Y131_CO6;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D = CLBLM_R_X93Y131_SLICE_X147Y131_DO6;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_AMUX = CLBLM_R_X93Y131_SLICE_X147Y131_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_BMUX = CLBLM_R_X93Y131_SLICE_X147Y131_B5Q;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A = CLBLM_R_X93Y132_SLICE_X146Y132_AO6;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B = CLBLM_R_X93Y132_SLICE_X146Y132_BO6;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C = CLBLM_R_X93Y132_SLICE_X146Y132_CO6;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D = CLBLM_R_X93Y132_SLICE_X146Y132_DO6;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_AMUX = CLBLM_R_X93Y132_SLICE_X146Y132_A5Q;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A = CLBLM_R_X93Y132_SLICE_X147Y132_AO6;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B = CLBLM_R_X93Y132_SLICE_X147Y132_BO6;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C = CLBLM_R_X93Y132_SLICE_X147Y132_CO6;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D = CLBLM_R_X93Y132_SLICE_X147Y132_DO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A = CLBLM_R_X93Y133_SLICE_X146Y133_AO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B = CLBLM_R_X93Y133_SLICE_X146Y133_BO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C = CLBLM_R_X93Y133_SLICE_X146Y133_CO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D = CLBLM_R_X93Y133_SLICE_X146Y133_DO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_AMUX = CLBLM_R_X93Y133_SLICE_X146Y133_A5Q;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_BMUX = CLBLM_R_X93Y133_SLICE_X146Y133_BO5;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_CMUX = CLBLM_R_X93Y133_SLICE_X146Y133_C5Q;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A = CLBLM_R_X93Y133_SLICE_X147Y133_AO6;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B = CLBLM_R_X93Y133_SLICE_X147Y133_BO6;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C = CLBLM_R_X93Y133_SLICE_X147Y133_CO6;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D = CLBLM_R_X93Y133_SLICE_X147Y133_DO6;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A = CLBLM_R_X95Y111_SLICE_X150Y111_AO6;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B = CLBLM_R_X95Y111_SLICE_X150Y111_BO6;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C = CLBLM_R_X95Y111_SLICE_X150Y111_CO6;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D = CLBLM_R_X95Y111_SLICE_X150Y111_DO6;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_AMUX = CLBLM_R_X95Y111_SLICE_X150Y111_A5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_BMUX = CLBLM_R_X95Y111_SLICE_X150Y111_B5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_CMUX = CLBLM_R_X95Y111_SLICE_X150Y111_C5Q;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A = CLBLM_R_X95Y111_SLICE_X151Y111_AO6;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B = CLBLM_R_X95Y111_SLICE_X151Y111_BO6;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C = CLBLM_R_X95Y111_SLICE_X151Y111_CO6;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D = CLBLM_R_X95Y111_SLICE_X151Y111_DO6;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_AMUX = CLBLM_R_X95Y111_SLICE_X151Y111_A5Q;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_BMUX = CLBLM_R_X95Y111_SLICE_X151Y111_B5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A = CLBLM_R_X95Y112_SLICE_X150Y112_AO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B = CLBLM_R_X95Y112_SLICE_X150Y112_BO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C = CLBLM_R_X95Y112_SLICE_X150Y112_CO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D = CLBLM_R_X95Y112_SLICE_X150Y112_DO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_AMUX = CLBLM_R_X95Y112_SLICE_X150Y112_A5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_BMUX = CLBLM_R_X95Y112_SLICE_X150Y112_B5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_CMUX = CLBLM_R_X95Y112_SLICE_X150Y112_CO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A = CLBLM_R_X95Y112_SLICE_X151Y112_AO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B = CLBLM_R_X95Y112_SLICE_X151Y112_BO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C = CLBLM_R_X95Y112_SLICE_X151Y112_CO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D = CLBLM_R_X95Y112_SLICE_X151Y112_DO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_AMUX = CLBLM_R_X95Y112_SLICE_X151Y112_AO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A = CLBLM_R_X95Y113_SLICE_X150Y113_AO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B = CLBLM_R_X95Y113_SLICE_X150Y113_BO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C = CLBLM_R_X95Y113_SLICE_X150Y113_CO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D = CLBLM_R_X95Y113_SLICE_X150Y113_DO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_AMUX = CLBLM_R_X95Y113_SLICE_X150Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_BMUX = CLBLM_R_X95Y113_SLICE_X150Y113_B5Q;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A = CLBLM_R_X95Y113_SLICE_X151Y113_AO6;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B = CLBLM_R_X95Y113_SLICE_X151Y113_BO6;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C = CLBLM_R_X95Y113_SLICE_X151Y113_CO6;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D = CLBLM_R_X95Y113_SLICE_X151Y113_DO6;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_AMUX = CLBLM_R_X95Y113_SLICE_X151Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_BMUX = CLBLM_R_X95Y113_SLICE_X151Y113_B5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A = CLBLM_R_X95Y114_SLICE_X150Y114_AO6;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B = CLBLM_R_X95Y114_SLICE_X150Y114_BO6;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C = CLBLM_R_X95Y114_SLICE_X150Y114_CO6;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D = CLBLM_R_X95Y114_SLICE_X150Y114_DO6;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_AMUX = CLBLM_R_X95Y114_SLICE_X150Y114_A5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_BMUX = CLBLM_R_X95Y114_SLICE_X150Y114_B5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_CMUX = CLBLM_R_X95Y114_SLICE_X150Y114_C5Q;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A = CLBLM_R_X95Y114_SLICE_X151Y114_AO6;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B = CLBLM_R_X95Y114_SLICE_X151Y114_BO6;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C = CLBLM_R_X95Y114_SLICE_X151Y114_CO6;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D = CLBLM_R_X95Y114_SLICE_X151Y114_DO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A = CLBLM_R_X95Y115_SLICE_X150Y115_AO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B = CLBLM_R_X95Y115_SLICE_X150Y115_BO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C = CLBLM_R_X95Y115_SLICE_X150Y115_CO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D = CLBLM_R_X95Y115_SLICE_X150Y115_DO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_AMUX = CLBLM_R_X95Y115_SLICE_X150Y115_A5Q;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_BMUX = CLBLM_R_X95Y115_SLICE_X150Y115_B5Q;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_CMUX = CLBLM_R_X95Y115_SLICE_X150Y115_C5Q;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_DMUX = CLBLM_R_X95Y115_SLICE_X150Y115_DO6;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A = CLBLM_R_X95Y115_SLICE_X151Y115_AO6;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B = CLBLM_R_X95Y115_SLICE_X151Y115_BO6;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C = CLBLM_R_X95Y115_SLICE_X151Y115_CO6;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D = CLBLM_R_X95Y115_SLICE_X151Y115_DO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A = CLBLM_R_X95Y116_SLICE_X150Y116_AO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B = CLBLM_R_X95Y116_SLICE_X150Y116_BO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C = CLBLM_R_X95Y116_SLICE_X150Y116_CO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D = CLBLM_R_X95Y116_SLICE_X150Y116_DO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_AMUX = CLBLM_R_X95Y116_SLICE_X150Y116_A5Q;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A = CLBLM_R_X95Y116_SLICE_X151Y116_AO6;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B = CLBLM_R_X95Y116_SLICE_X151Y116_BO6;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C = CLBLM_R_X95Y116_SLICE_X151Y116_CO6;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D = CLBLM_R_X95Y116_SLICE_X151Y116_DO6;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_AMUX = CLBLM_R_X95Y116_SLICE_X151Y116_A5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A = CLBLM_R_X95Y117_SLICE_X150Y117_AO6;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B = CLBLM_R_X95Y117_SLICE_X150Y117_BO6;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C = CLBLM_R_X95Y117_SLICE_X150Y117_CO6;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D = CLBLM_R_X95Y117_SLICE_X150Y117_DO6;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_AMUX = CLBLM_R_X95Y117_SLICE_X150Y117_A5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_BMUX = CLBLM_R_X95Y117_SLICE_X150Y117_B5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_CMUX = CLBLM_R_X95Y117_SLICE_X150Y117_C5Q;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A = CLBLM_R_X95Y117_SLICE_X151Y117_AO6;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B = CLBLM_R_X95Y117_SLICE_X151Y117_BO6;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C = CLBLM_R_X95Y117_SLICE_X151Y117_CO6;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D = CLBLM_R_X95Y117_SLICE_X151Y117_DO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A = CLBLM_R_X95Y118_SLICE_X150Y118_AO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B = CLBLM_R_X95Y118_SLICE_X150Y118_BO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C = CLBLM_R_X95Y118_SLICE_X150Y118_CO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D = CLBLM_R_X95Y118_SLICE_X150Y118_DO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_AMUX = CLBLM_R_X95Y118_SLICE_X150Y118_A5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_BMUX = CLBLM_R_X95Y118_SLICE_X150Y118_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_CMUX = CLBLM_R_X95Y118_SLICE_X150Y118_C5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_DMUX = CLBLM_R_X95Y118_SLICE_X150Y118_DO6;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A = CLBLM_R_X95Y118_SLICE_X151Y118_AO6;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B = CLBLM_R_X95Y118_SLICE_X151Y118_BO6;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C = CLBLM_R_X95Y118_SLICE_X151Y118_CO6;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D = CLBLM_R_X95Y118_SLICE_X151Y118_DO6;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_AMUX = CLBLM_R_X95Y118_SLICE_X151Y118_A5Q;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_BMUX = CLBLM_R_X95Y118_SLICE_X151Y118_B5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A = CLBLM_R_X95Y119_SLICE_X150Y119_AO6;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B = CLBLM_R_X95Y119_SLICE_X150Y119_BO6;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C = CLBLM_R_X95Y119_SLICE_X150Y119_CO6;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D = CLBLM_R_X95Y119_SLICE_X150Y119_DO6;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_AMUX = CLBLM_R_X95Y119_SLICE_X150Y119_A5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_BMUX = CLBLM_R_X95Y119_SLICE_X150Y119_B5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_CMUX = CLBLM_R_X95Y119_SLICE_X150Y119_C5Q;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A = CLBLM_R_X95Y119_SLICE_X151Y119_AO6;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B = CLBLM_R_X95Y119_SLICE_X151Y119_BO6;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C = CLBLM_R_X95Y119_SLICE_X151Y119_CO6;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D = CLBLM_R_X95Y119_SLICE_X151Y119_DO6;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A = CLBLM_R_X95Y120_SLICE_X150Y120_AO6;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B = CLBLM_R_X95Y120_SLICE_X150Y120_BO6;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C = CLBLM_R_X95Y120_SLICE_X150Y120_CO6;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D = CLBLM_R_X95Y120_SLICE_X150Y120_DO6;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_AMUX = CLBLM_R_X95Y120_SLICE_X150Y120_A5Q;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_BMUX = CLBLM_R_X95Y120_SLICE_X150Y120_B5Q;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A = CLBLM_R_X95Y120_SLICE_X151Y120_AO6;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B = CLBLM_R_X95Y120_SLICE_X151Y120_BO6;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C = CLBLM_R_X95Y120_SLICE_X151Y120_CO6;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D = CLBLM_R_X95Y120_SLICE_X151Y120_DO6;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_AMUX = CLBLM_R_X95Y120_SLICE_X151Y120_A5Q;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_BMUX = CLBLM_R_X95Y120_SLICE_X151Y120_B5Q;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A = CLBLM_R_X95Y121_SLICE_X150Y121_AO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B = CLBLM_R_X95Y121_SLICE_X150Y121_BO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C = CLBLM_R_X95Y121_SLICE_X150Y121_CO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D = CLBLM_R_X95Y121_SLICE_X150Y121_DO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_AMUX = CLBLM_R_X95Y121_SLICE_X150Y121_A5Q;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A = CLBLM_R_X95Y121_SLICE_X151Y121_AO6;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B = CLBLM_R_X95Y121_SLICE_X151Y121_BO6;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C = CLBLM_R_X95Y121_SLICE_X151Y121_CO6;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D = CLBLM_R_X95Y121_SLICE_X151Y121_DO6;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_AMUX = CLBLM_R_X95Y121_SLICE_X151Y121_A5Q;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_BMUX = CLBLM_R_X95Y121_SLICE_X151Y121_B5Q;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_CMUX = CLBLM_R_X95Y121_SLICE_X151Y121_CO6;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A = CLBLM_R_X95Y122_SLICE_X150Y122_AO6;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B = CLBLM_R_X95Y122_SLICE_X150Y122_BO6;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C = CLBLM_R_X95Y122_SLICE_X150Y122_CO6;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D = CLBLM_R_X95Y122_SLICE_X150Y122_DO6;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_AMUX = CLBLM_R_X95Y122_SLICE_X150Y122_A5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_BMUX = CLBLM_R_X95Y122_SLICE_X150Y122_B5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_CMUX = CLBLM_R_X95Y122_SLICE_X150Y122_C5Q;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A = CLBLM_R_X95Y122_SLICE_X151Y122_AO6;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B = CLBLM_R_X95Y122_SLICE_X151Y122_BO6;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C = CLBLM_R_X95Y122_SLICE_X151Y122_CO6;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D = CLBLM_R_X95Y122_SLICE_X151Y122_DO6;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A = CLBLM_R_X95Y123_SLICE_X150Y123_AO6;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B = CLBLM_R_X95Y123_SLICE_X150Y123_BO6;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C = CLBLM_R_X95Y123_SLICE_X150Y123_CO6;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D = CLBLM_R_X95Y123_SLICE_X150Y123_DO6;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_AMUX = CLBLM_R_X95Y123_SLICE_X150Y123_A5Q;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_BMUX = CLBLM_R_X95Y123_SLICE_X150Y123_B5Q;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A = CLBLM_R_X95Y123_SLICE_X151Y123_AO6;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B = CLBLM_R_X95Y123_SLICE_X151Y123_BO6;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C = CLBLM_R_X95Y123_SLICE_X151Y123_CO6;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D = CLBLM_R_X95Y123_SLICE_X151Y123_DO6;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_AMUX = CLBLM_R_X95Y123_SLICE_X151Y123_A5Q;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_BMUX = CLBLM_R_X95Y123_SLICE_X151Y123_B5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A = CLBLM_R_X95Y124_SLICE_X150Y124_AO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B = CLBLM_R_X95Y124_SLICE_X150Y124_BO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C = CLBLM_R_X95Y124_SLICE_X150Y124_CO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D = CLBLM_R_X95Y124_SLICE_X150Y124_DO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_AMUX = CLBLM_R_X95Y124_SLICE_X150Y124_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_BMUX = CLBLM_R_X95Y124_SLICE_X150Y124_B5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_CMUX = CLBLM_R_X95Y124_SLICE_X150Y124_C5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A = CLBLM_R_X95Y124_SLICE_X151Y124_AO6;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B = CLBLM_R_X95Y124_SLICE_X151Y124_BO6;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C = CLBLM_R_X95Y124_SLICE_X151Y124_CO6;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D = CLBLM_R_X95Y124_SLICE_X151Y124_DO6;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_AMUX = CLBLM_R_X95Y124_SLICE_X151Y124_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_BMUX = CLBLM_R_X95Y124_SLICE_X151Y124_BO5;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_CMUX = CLBLM_R_X95Y124_SLICE_X151Y124_C5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A = CLBLM_R_X95Y125_SLICE_X150Y125_AO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B = CLBLM_R_X95Y125_SLICE_X150Y125_BO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C = CLBLM_R_X95Y125_SLICE_X150Y125_CO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D = CLBLM_R_X95Y125_SLICE_X150Y125_DO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_AMUX = CLBLM_R_X95Y125_SLICE_X150Y125_A5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_BMUX = CLBLM_R_X95Y125_SLICE_X150Y125_B5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_CMUX = CLBLM_R_X95Y125_SLICE_X150Y125_CO5;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A = CLBLM_R_X95Y125_SLICE_X151Y125_AO6;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B = CLBLM_R_X95Y125_SLICE_X151Y125_BO6;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C = CLBLM_R_X95Y125_SLICE_X151Y125_CO6;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D = CLBLM_R_X95Y125_SLICE_X151Y125_DO6;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_AMUX = CLBLM_R_X95Y125_SLICE_X151Y125_A5Q;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A = CLBLM_R_X95Y126_SLICE_X150Y126_AO6;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B = CLBLM_R_X95Y126_SLICE_X150Y126_BO6;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C = CLBLM_R_X95Y126_SLICE_X150Y126_CO6;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D = CLBLM_R_X95Y126_SLICE_X150Y126_DO6;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_AMUX = CLBLM_R_X95Y126_SLICE_X150Y126_A5Q;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_BMUX = CLBLM_R_X95Y126_SLICE_X150Y126_B5Q;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A = CLBLM_R_X95Y126_SLICE_X151Y126_AO6;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B = CLBLM_R_X95Y126_SLICE_X151Y126_BO6;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C = CLBLM_R_X95Y126_SLICE_X151Y126_CO6;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D = CLBLM_R_X95Y126_SLICE_X151Y126_DO6;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_AMUX = CLBLM_R_X95Y126_SLICE_X151Y126_A5Q;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A = CLBLM_R_X95Y128_SLICE_X150Y128_AO6;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B = CLBLM_R_X95Y128_SLICE_X150Y128_BO6;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C = CLBLM_R_X95Y128_SLICE_X150Y128_CO6;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D = CLBLM_R_X95Y128_SLICE_X150Y128_DO6;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_BMUX = CLBLM_R_X95Y128_SLICE_X150Y128_B5Q;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A = CLBLM_R_X95Y128_SLICE_X151Y128_AO6;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B = CLBLM_R_X95Y128_SLICE_X151Y128_BO6;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C = CLBLM_R_X95Y128_SLICE_X151Y128_CO6;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D = CLBLM_R_X95Y128_SLICE_X151Y128_DO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A = CLBLM_R_X95Y129_SLICE_X150Y129_AO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B = CLBLM_R_X95Y129_SLICE_X150Y129_BO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C = CLBLM_R_X95Y129_SLICE_X150Y129_CO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D = CLBLM_R_X95Y129_SLICE_X150Y129_DO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_AMUX = CLBLM_R_X95Y129_SLICE_X150Y129_A5Q;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_BMUX = CLBLM_R_X95Y129_SLICE_X150Y129_BO5;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_CMUX = CLBLM_R_X95Y129_SLICE_X150Y129_C5Q;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A = CLBLM_R_X95Y129_SLICE_X151Y129_AO6;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B = CLBLM_R_X95Y129_SLICE_X151Y129_BO6;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C = CLBLM_R_X95Y129_SLICE_X151Y129_CO6;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D = CLBLM_R_X95Y129_SLICE_X151Y129_DO6;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_AMUX = CLBLM_R_X95Y129_SLICE_X151Y129_A5Q;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_BMUX = CLBLM_R_X95Y129_SLICE_X151Y129_B5Q;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_CMUX = CLBLM_R_X95Y129_SLICE_X151Y129_CO5;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_DMUX = CLBLM_R_X95Y129_SLICE_X151Y129_D5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A = CLBLM_R_X95Y130_SLICE_X150Y130_AO6;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B = CLBLM_R_X95Y130_SLICE_X150Y130_BO6;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C = CLBLM_R_X95Y130_SLICE_X150Y130_CO6;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D = CLBLM_R_X95Y130_SLICE_X150Y130_DO6;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_AMUX = CLBLM_R_X95Y130_SLICE_X150Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_BMUX = CLBLM_R_X95Y130_SLICE_X150Y130_BO5;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_CMUX = CLBLM_R_X95Y130_SLICE_X150Y130_C5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_DMUX = CLBLM_R_X95Y130_SLICE_X150Y130_DO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A = CLBLM_R_X95Y130_SLICE_X151Y130_AO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B = CLBLM_R_X95Y130_SLICE_X151Y130_BO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C = CLBLM_R_X95Y130_SLICE_X151Y130_CO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D = CLBLM_R_X95Y130_SLICE_X151Y130_DO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_AMUX = CLBLM_R_X95Y130_SLICE_X151Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_BMUX = CLBLM_R_X95Y130_SLICE_X151Y130_BO5;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_CMUX = CLBLM_R_X95Y130_SLICE_X151Y130_C5Q;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A = CLBLM_R_X95Y131_SLICE_X150Y131_AO6;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B = CLBLM_R_X95Y131_SLICE_X150Y131_BO6;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C = CLBLM_R_X95Y131_SLICE_X150Y131_CO6;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D = CLBLM_R_X95Y131_SLICE_X150Y131_DO6;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_AMUX = CLBLM_R_X95Y131_SLICE_X150Y131_A5Q;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_BMUX = CLBLM_R_X95Y131_SLICE_X150Y131_B5Q;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A = CLBLM_R_X95Y131_SLICE_X151Y131_AO6;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B = CLBLM_R_X95Y131_SLICE_X151Y131_BO6;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C = CLBLM_R_X95Y131_SLICE_X151Y131_CO6;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D = CLBLM_R_X95Y131_SLICE_X151Y131_DO6;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_AMUX = CLBLM_R_X95Y131_SLICE_X151Y131_A5Q;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_BMUX = CLBLM_R_X95Y131_SLICE_X151Y131_BO5;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_CMUX = CLBLM_R_X95Y131_SLICE_X151Y131_C5Q;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_DMUX = CLBLM_R_X95Y131_SLICE_X151Y131_D5Q;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A = CLBLM_R_X95Y132_SLICE_X150Y132_AO6;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B = CLBLM_R_X95Y132_SLICE_X150Y132_BO6;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C = CLBLM_R_X95Y132_SLICE_X150Y132_CO6;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D = CLBLM_R_X95Y132_SLICE_X150Y132_DO6;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_BMUX = CLBLM_R_X95Y132_SLICE_X150Y132_B5Q;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_CMUX = CLBLM_R_X95Y132_SLICE_X150Y132_C5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A = CLBLM_R_X95Y132_SLICE_X151Y132_AO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B = CLBLM_R_X95Y132_SLICE_X151Y132_BO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C = CLBLM_R_X95Y132_SLICE_X151Y132_CO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D = CLBLM_R_X95Y132_SLICE_X151Y132_DO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_AMUX = CLBLM_R_X95Y132_SLICE_X151Y132_A5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_BMUX = CLBLM_R_X95Y132_SLICE_X151Y132_B5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_DMUX = CLBLM_R_X95Y132_SLICE_X151Y132_DO5;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A = CLBLM_R_X97Y111_SLICE_X152Y111_AO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B = CLBLM_R_X97Y111_SLICE_X152Y111_BO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C = CLBLM_R_X97Y111_SLICE_X152Y111_CO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D = CLBLM_R_X97Y111_SLICE_X152Y111_DO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_AMUX = CLBLM_R_X97Y111_SLICE_X152Y111_A5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_BMUX = CLBLM_R_X97Y111_SLICE_X152Y111_B5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_CMUX = CLBLM_R_X97Y111_SLICE_X152Y111_CO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A = CLBLM_R_X97Y111_SLICE_X153Y111_AO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B = CLBLM_R_X97Y111_SLICE_X153Y111_BO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C = CLBLM_R_X97Y111_SLICE_X153Y111_CO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D = CLBLM_R_X97Y111_SLICE_X153Y111_DO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_AMUX = CLBLM_R_X97Y111_SLICE_X153Y111_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A = CLBLM_R_X97Y112_SLICE_X152Y112_AO6;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B = CLBLM_R_X97Y112_SLICE_X152Y112_BO6;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C = CLBLM_R_X97Y112_SLICE_X152Y112_CO6;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D = CLBLM_R_X97Y112_SLICE_X152Y112_DO6;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_AMUX = CLBLM_R_X97Y112_SLICE_X152Y112_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_BMUX = CLBLM_R_X97Y112_SLICE_X152Y112_B5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_CMUX = CLBLM_R_X97Y112_SLICE_X152Y112_C5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A = CLBLM_R_X97Y112_SLICE_X153Y112_AO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B = CLBLM_R_X97Y112_SLICE_X153Y112_BO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C = CLBLM_R_X97Y112_SLICE_X153Y112_CO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D = CLBLM_R_X97Y112_SLICE_X153Y112_DO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_AMUX = CLBLM_R_X97Y112_SLICE_X153Y112_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_BMUX = CLBLM_R_X97Y112_SLICE_X153Y112_B5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_CMUX = CLBLM_R_X97Y112_SLICE_X153Y112_CO6;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A = CLBLM_R_X97Y113_SLICE_X152Y113_AO6;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B = CLBLM_R_X97Y113_SLICE_X152Y113_BO6;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C = CLBLM_R_X97Y113_SLICE_X152Y113_CO6;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D = CLBLM_R_X97Y113_SLICE_X152Y113_DO6;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_AMUX = CLBLM_R_X97Y113_SLICE_X152Y113_A5Q;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A = CLBLM_R_X97Y113_SLICE_X153Y113_AO6;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B = CLBLM_R_X97Y113_SLICE_X153Y113_BO6;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C = CLBLM_R_X97Y113_SLICE_X153Y113_CO6;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D = CLBLM_R_X97Y113_SLICE_X153Y113_DO6;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A = CLBLM_R_X97Y115_SLICE_X152Y115_AO6;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B = CLBLM_R_X97Y115_SLICE_X152Y115_BO6;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C = CLBLM_R_X97Y115_SLICE_X152Y115_CO6;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D = CLBLM_R_X97Y115_SLICE_X152Y115_DO6;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_AMUX = CLBLM_R_X97Y115_SLICE_X152Y115_A5Q;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A = CLBLM_R_X97Y115_SLICE_X153Y115_AO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B = CLBLM_R_X97Y115_SLICE_X153Y115_BO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C = CLBLM_R_X97Y115_SLICE_X153Y115_CO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D = CLBLM_R_X97Y115_SLICE_X153Y115_DO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_AMUX = CLBLM_R_X97Y115_SLICE_X153Y115_A5Q;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_BMUX = CLBLM_R_X97Y115_SLICE_X153Y115_B5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A = CLBLM_R_X97Y116_SLICE_X152Y116_AO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B = CLBLM_R_X97Y116_SLICE_X152Y116_BO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C = CLBLM_R_X97Y116_SLICE_X152Y116_CO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D = CLBLM_R_X97Y116_SLICE_X152Y116_DO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_AMUX = CLBLM_R_X97Y116_SLICE_X152Y116_A5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_BMUX = CLBLM_R_X97Y116_SLICE_X152Y116_B5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_CMUX = CLBLM_R_X97Y116_SLICE_X152Y116_CO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A = CLBLM_R_X97Y116_SLICE_X153Y116_AO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B = CLBLM_R_X97Y116_SLICE_X153Y116_BO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C = CLBLM_R_X97Y116_SLICE_X153Y116_CO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D = CLBLM_R_X97Y116_SLICE_X153Y116_DO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_AMUX = CLBLM_R_X97Y116_SLICE_X153Y116_A5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_BMUX = CLBLM_R_X97Y116_SLICE_X153Y116_B5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_CMUX = CLBLM_R_X97Y116_SLICE_X153Y116_C5Q;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A = CLBLM_R_X97Y117_SLICE_X152Y117_AO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B = CLBLM_R_X97Y117_SLICE_X152Y117_BO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C = CLBLM_R_X97Y117_SLICE_X152Y117_CO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D = CLBLM_R_X97Y117_SLICE_X152Y117_DO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_AMUX = CLBLM_R_X97Y117_SLICE_X152Y117_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_BMUX = CLBLM_R_X97Y117_SLICE_X152Y117_B5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A = CLBLM_R_X97Y117_SLICE_X153Y117_AO6;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B = CLBLM_R_X97Y117_SLICE_X153Y117_BO6;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C = CLBLM_R_X97Y117_SLICE_X153Y117_CO6;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D = CLBLM_R_X97Y117_SLICE_X153Y117_DO6;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_AMUX = CLBLM_R_X97Y117_SLICE_X153Y117_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_CMUX = CLBLM_R_X97Y117_SLICE_X153Y117_C5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_DMUX = CLBLM_R_X97Y117_SLICE_X153Y117_DO5;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A = CLBLM_R_X97Y118_SLICE_X152Y118_AO6;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B = CLBLM_R_X97Y118_SLICE_X152Y118_BO6;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C = CLBLM_R_X97Y118_SLICE_X152Y118_CO6;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D = CLBLM_R_X97Y118_SLICE_X152Y118_DO6;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_AMUX = CLBLM_R_X97Y118_SLICE_X152Y118_A5Q;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_BMUX = CLBLM_R_X97Y118_SLICE_X152Y118_BO5;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_CMUX = CLBLM_R_X97Y118_SLICE_X152Y118_C5Q;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A = CLBLM_R_X97Y118_SLICE_X153Y118_AO6;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B = CLBLM_R_X97Y118_SLICE_X153Y118_BO6;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C = CLBLM_R_X97Y118_SLICE_X153Y118_CO6;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D = CLBLM_R_X97Y118_SLICE_X153Y118_DO6;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_BMUX = CLBLM_R_X97Y118_SLICE_X153Y118_B5Q;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_CMUX = CLBLM_R_X97Y118_SLICE_X153Y118_C5Q;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A = CLBLM_R_X97Y119_SLICE_X152Y119_AO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B = CLBLM_R_X97Y119_SLICE_X152Y119_BO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C = CLBLM_R_X97Y119_SLICE_X152Y119_CO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D = CLBLM_R_X97Y119_SLICE_X152Y119_DO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_AMUX = CLBLM_R_X97Y119_SLICE_X152Y119_A5Q;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_BMUX = CLBLM_R_X97Y119_SLICE_X152Y119_B5Q;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A = CLBLM_R_X97Y119_SLICE_X153Y119_AO6;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B = CLBLM_R_X97Y119_SLICE_X153Y119_BO6;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C = CLBLM_R_X97Y119_SLICE_X153Y119_CO6;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D = CLBLM_R_X97Y119_SLICE_X153Y119_DO6;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_AMUX = CLBLM_R_X97Y119_SLICE_X153Y119_A5Q;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_CMUX = CLBLM_R_X97Y119_SLICE_X153Y119_C5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A = CLBLM_R_X97Y120_SLICE_X152Y120_AO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B = CLBLM_R_X97Y120_SLICE_X152Y120_BO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C = CLBLM_R_X97Y120_SLICE_X152Y120_CO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D = CLBLM_R_X97Y120_SLICE_X152Y120_DO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_AMUX = CLBLM_R_X97Y120_SLICE_X152Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_CMUX = CLBLM_R_X97Y120_SLICE_X152Y120_CO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A = CLBLM_R_X97Y120_SLICE_X153Y120_AO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B = CLBLM_R_X97Y120_SLICE_X153Y120_BO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C = CLBLM_R_X97Y120_SLICE_X153Y120_CO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D = CLBLM_R_X97Y120_SLICE_X153Y120_DO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_AMUX = CLBLM_R_X97Y120_SLICE_X153Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_BMUX = CLBLM_R_X97Y120_SLICE_X153Y120_B5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_CMUX = CLBLM_R_X97Y120_SLICE_X153Y120_C5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_DMUX = CLBLM_R_X97Y120_SLICE_X153Y120_D5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A = CLBLM_R_X97Y121_SLICE_X152Y121_AO6;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B = CLBLM_R_X97Y121_SLICE_X152Y121_BO6;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C = CLBLM_R_X97Y121_SLICE_X152Y121_CO6;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D = CLBLM_R_X97Y121_SLICE_X152Y121_DO6;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_AMUX = CLBLM_R_X97Y121_SLICE_X152Y121_A5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_BMUX = CLBLM_R_X97Y121_SLICE_X152Y121_B5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_CMUX = CLBLM_R_X97Y121_SLICE_X152Y121_C5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A = CLBLM_R_X97Y121_SLICE_X153Y121_AO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B = CLBLM_R_X97Y121_SLICE_X153Y121_BO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C = CLBLM_R_X97Y121_SLICE_X153Y121_CO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D = CLBLM_R_X97Y121_SLICE_X153Y121_DO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_AMUX = CLBLM_R_X97Y121_SLICE_X153Y121_A5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_BMUX = CLBLM_R_X97Y121_SLICE_X153Y121_B5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_CMUX = CLBLM_R_X97Y121_SLICE_X153Y121_C5Q;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A = CLBLM_R_X97Y122_SLICE_X152Y122_AO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B = CLBLM_R_X97Y122_SLICE_X152Y122_BO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C = CLBLM_R_X97Y122_SLICE_X152Y122_CO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D = CLBLM_R_X97Y122_SLICE_X152Y122_DO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_AMUX = CLBLM_R_X97Y122_SLICE_X152Y122_A5Q;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_DMUX = CLBLM_R_X97Y122_SLICE_X152Y122_D5Q;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A = CLBLM_R_X97Y122_SLICE_X153Y122_AO6;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B = CLBLM_R_X97Y122_SLICE_X153Y122_BO6;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C = CLBLM_R_X97Y122_SLICE_X153Y122_CO6;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D = CLBLM_R_X97Y122_SLICE_X153Y122_DO6;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_BMUX = CLBLM_R_X97Y122_SLICE_X153Y122_B5Q;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_CMUX = CLBLM_R_X97Y122_SLICE_X153Y122_C5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A = CLBLM_R_X97Y123_SLICE_X152Y123_AO6;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B = CLBLM_R_X97Y123_SLICE_X152Y123_BO6;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C = CLBLM_R_X97Y123_SLICE_X152Y123_CO6;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D = CLBLM_R_X97Y123_SLICE_X152Y123_DO6;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_AMUX = CLBLM_R_X97Y123_SLICE_X152Y123_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_BMUX = CLBLM_R_X97Y123_SLICE_X152Y123_B5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_CMUX = CLBLM_R_X97Y123_SLICE_X152Y123_C5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A = CLBLM_R_X97Y123_SLICE_X153Y123_AO6;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B = CLBLM_R_X97Y123_SLICE_X153Y123_BO6;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C = CLBLM_R_X97Y123_SLICE_X153Y123_CO6;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D = CLBLM_R_X97Y123_SLICE_X153Y123_DO6;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_AMUX = CLBLM_R_X97Y123_SLICE_X153Y123_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_BMUX = CLBLM_R_X97Y123_SLICE_X153Y123_B5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_CMUX = CLBLM_R_X97Y123_SLICE_X153Y123_C5Q;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A = CLBLM_R_X97Y124_SLICE_X152Y124_AO6;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B = CLBLM_R_X97Y124_SLICE_X152Y124_BO6;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C = CLBLM_R_X97Y124_SLICE_X152Y124_CO6;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D = CLBLM_R_X97Y124_SLICE_X152Y124_DO6;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_AMUX = CLBLM_R_X97Y124_SLICE_X152Y124_A5Q;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_BMUX = CLBLM_R_X97Y124_SLICE_X152Y124_B5Q;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A = CLBLM_R_X97Y124_SLICE_X153Y124_AO6;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B = CLBLM_R_X97Y124_SLICE_X153Y124_BO6;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C = CLBLM_R_X97Y124_SLICE_X153Y124_CO6;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D = CLBLM_R_X97Y124_SLICE_X153Y124_DO6;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A = CLBLM_R_X97Y125_SLICE_X152Y125_AO6;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B = CLBLM_R_X97Y125_SLICE_X152Y125_BO6;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C = CLBLM_R_X97Y125_SLICE_X152Y125_CO6;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D = CLBLM_R_X97Y125_SLICE_X152Y125_DO6;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_AMUX = CLBLM_R_X97Y125_SLICE_X152Y125_A5Q;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_BMUX = CLBLM_R_X97Y125_SLICE_X152Y125_B5Q;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A = CLBLM_R_X97Y125_SLICE_X153Y125_AO6;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B = CLBLM_R_X97Y125_SLICE_X153Y125_BO6;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C = CLBLM_R_X97Y125_SLICE_X153Y125_CO6;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D = CLBLM_R_X97Y125_SLICE_X153Y125_DO6;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_AMUX = CLBLM_R_X97Y125_SLICE_X153Y125_A5Q;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_BMUX = CLBLM_R_X97Y125_SLICE_X153Y125_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A = CLBLM_R_X97Y126_SLICE_X152Y126_AO6;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B = CLBLM_R_X97Y126_SLICE_X152Y126_BO6;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C = CLBLM_R_X97Y126_SLICE_X152Y126_CO6;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D = CLBLM_R_X97Y126_SLICE_X152Y126_DO6;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_AMUX = CLBLM_R_X97Y126_SLICE_X152Y126_A5Q;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_BMUX = CLBLM_R_X97Y126_SLICE_X152Y126_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A = CLBLM_R_X97Y126_SLICE_X153Y126_AO6;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B = CLBLM_R_X97Y126_SLICE_X153Y126_BO6;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C = CLBLM_R_X97Y126_SLICE_X153Y126_CO6;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D = CLBLM_R_X97Y126_SLICE_X153Y126_DO6;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_BMUX = CLBLM_R_X97Y126_SLICE_X153Y126_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_CMUX = CLBLM_R_X97Y126_SLICE_X153Y126_C5Q;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A = CLBLM_R_X97Y127_SLICE_X152Y127_AO6;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B = CLBLM_R_X97Y127_SLICE_X152Y127_BO6;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C = CLBLM_R_X97Y127_SLICE_X152Y127_CO6;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D = CLBLM_R_X97Y127_SLICE_X152Y127_DO6;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_AMUX = CLBLM_R_X97Y127_SLICE_X152Y127_A5Q;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_BMUX = CLBLM_R_X97Y127_SLICE_X152Y127_B5Q;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_CMUX = CLBLM_R_X97Y127_SLICE_X152Y127_CO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A = CLBLM_R_X97Y127_SLICE_X153Y127_AO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B = CLBLM_R_X97Y127_SLICE_X153Y127_BO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C = CLBLM_R_X97Y127_SLICE_X153Y127_CO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D = CLBLM_R_X97Y127_SLICE_X153Y127_DO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_AMUX = CLBLM_R_X97Y127_SLICE_X153Y127_A5Q;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A = CLBLM_R_X97Y128_SLICE_X152Y128_AO6;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B = CLBLM_R_X97Y128_SLICE_X152Y128_BO6;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C = CLBLM_R_X97Y128_SLICE_X152Y128_CO6;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D = CLBLM_R_X97Y128_SLICE_X152Y128_DO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A = CLBLM_R_X97Y128_SLICE_X153Y128_AO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B = CLBLM_R_X97Y128_SLICE_X153Y128_BO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C = CLBLM_R_X97Y128_SLICE_X153Y128_CO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D = CLBLM_R_X97Y128_SLICE_X153Y128_DO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_AMUX = CLBLM_R_X97Y128_SLICE_X153Y128_A5Q;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_BMUX = CLBLM_R_X97Y128_SLICE_X153Y128_BO5;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_CMUX = CLBLM_R_X97Y128_SLICE_X153Y128_C5Q;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A = CLBLM_R_X97Y129_SLICE_X152Y129_AO6;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B = CLBLM_R_X97Y129_SLICE_X152Y129_BO6;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C = CLBLM_R_X97Y129_SLICE_X152Y129_CO6;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D = CLBLM_R_X97Y129_SLICE_X152Y129_DO6;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_AMUX = CLBLM_R_X97Y129_SLICE_X152Y129_A5Q;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_BMUX = CLBLM_R_X97Y129_SLICE_X152Y129_B5Q;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A = CLBLM_R_X97Y129_SLICE_X153Y129_AO6;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B = CLBLM_R_X97Y129_SLICE_X153Y129_BO6;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C = CLBLM_R_X97Y129_SLICE_X153Y129_CO6;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D = CLBLM_R_X97Y129_SLICE_X153Y129_DO6;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A = CLBLM_R_X97Y130_SLICE_X152Y130_AO6;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B = CLBLM_R_X97Y130_SLICE_X152Y130_BO6;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C = CLBLM_R_X97Y130_SLICE_X152Y130_CO6;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D = CLBLM_R_X97Y130_SLICE_X152Y130_DO6;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_BMUX = CLBLM_R_X97Y130_SLICE_X152Y130_B5Q;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A = CLBLM_R_X97Y130_SLICE_X153Y130_AO6;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B = CLBLM_R_X97Y130_SLICE_X153Y130_BO6;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C = CLBLM_R_X97Y130_SLICE_X153Y130_CO6;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D = CLBLM_R_X97Y130_SLICE_X153Y130_DO6;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_AMUX = CLBLM_R_X97Y130_SLICE_X153Y130_A5Q;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A = CLBLM_R_X97Y131_SLICE_X152Y131_AO6;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B = CLBLM_R_X97Y131_SLICE_X152Y131_BO6;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C = CLBLM_R_X97Y131_SLICE_X152Y131_CO6;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D = CLBLM_R_X97Y131_SLICE_X152Y131_DO6;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_BMUX = CLBLM_R_X97Y131_SLICE_X152Y131_B5Q;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A = CLBLM_R_X97Y131_SLICE_X153Y131_AO6;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B = CLBLM_R_X97Y131_SLICE_X153Y131_BO6;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C = CLBLM_R_X97Y131_SLICE_X153Y131_CO6;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D = CLBLM_R_X97Y131_SLICE_X153Y131_DO6;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_BMUX = CLBLM_R_X97Y131_SLICE_X153Y131_B5Q;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_CMUX = CLBLM_R_X97Y131_SLICE_X153Y131_C5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A = CLBLM_R_X97Y132_SLICE_X152Y132_AO6;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B = CLBLM_R_X97Y132_SLICE_X152Y132_BO6;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C = CLBLM_R_X97Y132_SLICE_X152Y132_CO6;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D = CLBLM_R_X97Y132_SLICE_X152Y132_DO6;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_AMUX = CLBLM_R_X97Y132_SLICE_X152Y132_A5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_BMUX = CLBLM_R_X97Y132_SLICE_X152Y132_B5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_CMUX = CLBLM_R_X97Y132_SLICE_X152Y132_CO5;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_DMUX = CLBLM_R_X97Y132_SLICE_X152Y132_D5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A = CLBLM_R_X97Y132_SLICE_X153Y132_AO6;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B = CLBLM_R_X97Y132_SLICE_X153Y132_BO6;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C = CLBLM_R_X97Y132_SLICE_X153Y132_CO6;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D = CLBLM_R_X97Y132_SLICE_X153Y132_DO6;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_AMUX = CLBLM_R_X97Y132_SLICE_X153Y132_A5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_BMUX = CLBLM_R_X97Y132_SLICE_X153Y132_B5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_CMUX = CLBLM_R_X97Y132_SLICE_X153Y132_C5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_DMUX = CLBLM_R_X97Y132_SLICE_X153Y132_DO6;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A = CLBLM_R_X97Y133_SLICE_X152Y133_AO6;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B = CLBLM_R_X97Y133_SLICE_X152Y133_BO6;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C = CLBLM_R_X97Y133_SLICE_X152Y133_CO6;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D = CLBLM_R_X97Y133_SLICE_X152Y133_DO6;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_AMUX = CLBLM_R_X97Y133_SLICE_X152Y133_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_BMUX = CLBLM_R_X97Y133_SLICE_X152Y133_BO5;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_CMUX = CLBLM_R_X97Y133_SLICE_X152Y133_C5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A = CLBLM_R_X97Y133_SLICE_X153Y133_AO6;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B = CLBLM_R_X97Y133_SLICE_X153Y133_BO6;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C = CLBLM_R_X97Y133_SLICE_X153Y133_CO6;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D = CLBLM_R_X97Y133_SLICE_X153Y133_DO6;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_AMUX = CLBLM_R_X97Y133_SLICE_X153Y133_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_BMUX = CLBLM_R_X97Y133_SLICE_X153Y133_BO5;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_CMUX = CLBLM_R_X97Y133_SLICE_X153Y133_C5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_DMUX = CLBLM_R_X97Y133_SLICE_X153Y133_DO6;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A = CLBLM_R_X101Y110_SLICE_X158Y110_AO6;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B = CLBLM_R_X101Y110_SLICE_X158Y110_BO6;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C = CLBLM_R_X101Y110_SLICE_X158Y110_CO6;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D = CLBLM_R_X101Y110_SLICE_X158Y110_DO6;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_AMUX = CLBLM_R_X101Y110_SLICE_X158Y110_A5Q;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_BMUX = CLBLM_R_X101Y110_SLICE_X158Y110_B5Q;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A = CLBLM_R_X101Y110_SLICE_X159Y110_AO6;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B = CLBLM_R_X101Y110_SLICE_X159Y110_BO6;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C = CLBLM_R_X101Y110_SLICE_X159Y110_CO6;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D = CLBLM_R_X101Y110_SLICE_X159Y110_DO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A = CLBLM_R_X101Y111_SLICE_X158Y111_AO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B = CLBLM_R_X101Y111_SLICE_X158Y111_BO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C = CLBLM_R_X101Y111_SLICE_X158Y111_CO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D = CLBLM_R_X101Y111_SLICE_X158Y111_DO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_AMUX = CLBLM_R_X101Y111_SLICE_X158Y111_A5Q;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_BMUX = CLBLM_R_X101Y111_SLICE_X158Y111_B5Q;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_CMUX = CLBLM_R_X101Y111_SLICE_X158Y111_CO6;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A = CLBLM_R_X101Y111_SLICE_X159Y111_AO6;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B = CLBLM_R_X101Y111_SLICE_X159Y111_BO6;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C = CLBLM_R_X101Y111_SLICE_X159Y111_CO6;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D = CLBLM_R_X101Y111_SLICE_X159Y111_DO6;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_AMUX = CLBLM_R_X101Y111_SLICE_X159Y111_A5Q;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_BMUX = CLBLM_R_X101Y111_SLICE_X159Y111_B5Q;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A = CLBLM_R_X101Y112_SLICE_X158Y112_AO6;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B = CLBLM_R_X101Y112_SLICE_X158Y112_BO6;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C = CLBLM_R_X101Y112_SLICE_X158Y112_CO6;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D = CLBLM_R_X101Y112_SLICE_X158Y112_DO6;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_AMUX = CLBLM_R_X101Y112_SLICE_X158Y112_A5Q;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_BMUX = CLBLM_R_X101Y112_SLICE_X158Y112_B5Q;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A = CLBLM_R_X101Y112_SLICE_X159Y112_AO6;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B = CLBLM_R_X101Y112_SLICE_X159Y112_BO6;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C = CLBLM_R_X101Y112_SLICE_X159Y112_CO6;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D = CLBLM_R_X101Y112_SLICE_X159Y112_DO6;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_AMUX = CLBLM_R_X101Y112_SLICE_X159Y112_A5Q;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_BMUX = CLBLM_R_X101Y112_SLICE_X159Y112_B5Q;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_CMUX = CLBLM_R_X101Y112_SLICE_X159Y112_C5Q;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A = CLBLM_R_X101Y113_SLICE_X158Y113_AO6;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B = CLBLM_R_X101Y113_SLICE_X158Y113_BO6;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C = CLBLM_R_X101Y113_SLICE_X158Y113_CO6;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D = CLBLM_R_X101Y113_SLICE_X158Y113_DO6;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_AMUX = CLBLM_R_X101Y113_SLICE_X158Y113_A5Q;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_BMUX = CLBLM_R_X101Y113_SLICE_X158Y113_B5Q;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A = CLBLM_R_X101Y113_SLICE_X159Y113_AO6;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B = CLBLM_R_X101Y113_SLICE_X159Y113_BO6;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C = CLBLM_R_X101Y113_SLICE_X159Y113_CO6;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D = CLBLM_R_X101Y113_SLICE_X159Y113_DO6;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_AMUX = CLBLM_R_X101Y113_SLICE_X159Y113_AO5;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_BMUX = CLBLM_R_X101Y113_SLICE_X159Y113_BO5;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_CMUX = CLBLM_R_X101Y113_SLICE_X159Y113_C5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A = CLBLM_R_X101Y114_SLICE_X158Y114_AO6;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B = CLBLM_R_X101Y114_SLICE_X158Y114_BO6;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C = CLBLM_R_X101Y114_SLICE_X158Y114_CO6;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D = CLBLM_R_X101Y114_SLICE_X158Y114_DO6;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_AMUX = CLBLM_R_X101Y114_SLICE_X158Y114_A5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_BMUX = CLBLM_R_X101Y114_SLICE_X158Y114_B5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_CMUX = CLBLM_R_X101Y114_SLICE_X158Y114_CO6;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A = CLBLM_R_X101Y114_SLICE_X159Y114_AO6;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B = CLBLM_R_X101Y114_SLICE_X159Y114_BO6;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C = CLBLM_R_X101Y114_SLICE_X159Y114_CO6;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D = CLBLM_R_X101Y114_SLICE_X159Y114_DO6;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A = CLBLM_R_X101Y115_SLICE_X158Y115_AO6;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B = CLBLM_R_X101Y115_SLICE_X158Y115_BO6;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C = CLBLM_R_X101Y115_SLICE_X158Y115_CO6;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D = CLBLM_R_X101Y115_SLICE_X158Y115_DO6;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_AMUX = CLBLM_R_X101Y115_SLICE_X158Y115_A5Q;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_BMUX = CLBLM_R_X101Y115_SLICE_X158Y115_B5Q;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A = CLBLM_R_X101Y115_SLICE_X159Y115_AO6;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B = CLBLM_R_X101Y115_SLICE_X159Y115_BO6;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C = CLBLM_R_X101Y115_SLICE_X159Y115_CO6;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D = CLBLM_R_X101Y115_SLICE_X159Y115_DO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A = CLBLM_R_X101Y116_SLICE_X158Y116_AO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B = CLBLM_R_X101Y116_SLICE_X158Y116_BO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C = CLBLM_R_X101Y116_SLICE_X158Y116_CO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D = CLBLM_R_X101Y116_SLICE_X158Y116_DO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_AMUX = CLBLM_R_X101Y116_SLICE_X158Y116_A5Q;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_BMUX = CLBLM_R_X101Y116_SLICE_X158Y116_B5Q;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_CMUX = CLBLM_R_X101Y116_SLICE_X158Y116_CO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A = CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B = CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C = CLBLM_R_X101Y116_SLICE_X159Y116_CO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D = CLBLM_R_X101Y116_SLICE_X159Y116_DO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_AMUX = CLBLM_R_X101Y116_SLICE_X159Y116_AO5;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_BMUX = CLBLM_R_X101Y116_SLICE_X159Y116_BO5;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_CMUX = CLBLM_R_X101Y116_SLICE_X159Y116_C5Q;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A = CLBLM_R_X101Y117_SLICE_X158Y117_AO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B = CLBLM_R_X101Y117_SLICE_X158Y117_BO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C = CLBLM_R_X101Y117_SLICE_X158Y117_CO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D = CLBLM_R_X101Y117_SLICE_X158Y117_DO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_BMUX = CLBLM_R_X101Y117_SLICE_X158Y117_B5Q;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_CMUX = CLBLM_R_X101Y117_SLICE_X158Y117_CO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A = CLBLM_R_X101Y117_SLICE_X159Y117_AO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B = CLBLM_R_X101Y117_SLICE_X159Y117_BO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C = CLBLM_R_X101Y117_SLICE_X159Y117_CO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D = CLBLM_R_X101Y117_SLICE_X159Y117_DO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_AMUX = CLBLM_R_X101Y117_SLICE_X159Y117_AO5;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_BMUX = CLBLM_R_X101Y117_SLICE_X159Y117_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A = CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B = CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C = CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_AMUX = CLBLM_R_X101Y118_SLICE_X158Y118_A5Q;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_BMUX = CLBLM_R_X101Y118_SLICE_X158Y118_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A = CLBLM_R_X101Y118_SLICE_X159Y118_AO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B = CLBLM_R_X101Y118_SLICE_X159Y118_BO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C = CLBLM_R_X101Y118_SLICE_X159Y118_CO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D = CLBLM_R_X101Y118_SLICE_X159Y118_DO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_AMUX = CLBLM_R_X101Y118_SLICE_X159Y118_A5Q;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_BMUX = CLBLM_R_X101Y118_SLICE_X159Y118_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_CMUX = CLBLM_R_X101Y118_SLICE_X159Y118_CO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A = CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B = CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C = CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D = CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_AMUX = CLBLM_R_X101Y119_SLICE_X158Y119_A5Q;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A = CLBLM_R_X101Y119_SLICE_X159Y119_AO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B = CLBLM_R_X101Y119_SLICE_X159Y119_BO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C = CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D = CLBLM_R_X101Y119_SLICE_X159Y119_DO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_AMUX = CLBLM_R_X101Y119_SLICE_X159Y119_A5Q;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_BMUX = CLBLM_R_X101Y119_SLICE_X159Y119_B5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A = CLBLM_R_X101Y120_SLICE_X158Y120_AO6;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B = CLBLM_R_X101Y120_SLICE_X158Y120_BO6;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C = CLBLM_R_X101Y120_SLICE_X158Y120_CO6;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D = CLBLM_R_X101Y120_SLICE_X158Y120_DO6;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_AMUX = CLBLM_R_X101Y120_SLICE_X158Y120_A5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_BMUX = CLBLM_R_X101Y120_SLICE_X158Y120_BO5;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_CMUX = CLBLM_R_X101Y120_SLICE_X158Y120_C5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_DMUX = CLBLM_R_X101Y120_SLICE_X158Y120_DO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A = CLBLM_R_X101Y120_SLICE_X159Y120_AO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B = CLBLM_R_X101Y120_SLICE_X159Y120_BO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C = CLBLM_R_X101Y120_SLICE_X159Y120_CO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D = CLBLM_R_X101Y120_SLICE_X159Y120_DO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_BMUX = CLBLM_R_X101Y120_SLICE_X159Y120_B5Q;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A = CLBLM_R_X101Y121_SLICE_X158Y121_AO6;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B = CLBLM_R_X101Y121_SLICE_X158Y121_BO6;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C = CLBLM_R_X101Y121_SLICE_X158Y121_CO6;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D = CLBLM_R_X101Y121_SLICE_X158Y121_DO6;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_AMUX = CLBLM_R_X101Y121_SLICE_X158Y121_A5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A = CLBLM_R_X101Y121_SLICE_X159Y121_AO6;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B = CLBLM_R_X101Y121_SLICE_X159Y121_BO6;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C = CLBLM_R_X101Y121_SLICE_X159Y121_CO6;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D = CLBLM_R_X101Y121_SLICE_X159Y121_DO6;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_AMUX = CLBLM_R_X101Y121_SLICE_X159Y121_A5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_BMUX = CLBLM_R_X101Y121_SLICE_X159Y121_B5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_CMUX = CLBLM_R_X101Y121_SLICE_X159Y121_C5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_DMUX = CLBLM_R_X101Y121_SLICE_X159Y121_DO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A = CLBLM_R_X101Y122_SLICE_X158Y122_AO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B = CLBLM_R_X101Y122_SLICE_X158Y122_BO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C = CLBLM_R_X101Y122_SLICE_X158Y122_CO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D = CLBLM_R_X101Y122_SLICE_X158Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_AMUX = CLBLM_R_X101Y122_SLICE_X158Y122_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_BMUX = CLBLM_R_X101Y122_SLICE_X158Y122_B5Q;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_DMUX = CLBLM_R_X101Y122_SLICE_X158Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A = CLBLM_R_X101Y122_SLICE_X159Y122_AO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B = CLBLM_R_X101Y122_SLICE_X159Y122_BO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C = CLBLM_R_X101Y122_SLICE_X159Y122_CO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D = CLBLM_R_X101Y122_SLICE_X159Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_AMUX = CLBLM_R_X101Y122_SLICE_X159Y122_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_BMUX = CLBLM_R_X101Y122_SLICE_X159Y122_B5Q;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B = CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D = CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_AMUX = CLBLM_R_X101Y123_SLICE_X158Y123_A5Q;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_BMUX = CLBLM_R_X101Y123_SLICE_X158Y123_B5Q;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_DMUX = CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A = CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B = CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C = CLBLM_R_X101Y123_SLICE_X159Y123_CO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D = CLBLM_R_X101Y123_SLICE_X159Y123_DO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_AMUX = CLBLM_R_X101Y123_SLICE_X159Y123_A5Q;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_CMUX = CLBLM_R_X101Y123_SLICE_X159Y123_C5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A = CLBLM_R_X101Y124_SLICE_X158Y124_AO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B = CLBLM_R_X101Y124_SLICE_X158Y124_BO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_AMUX = CLBLM_R_X101Y124_SLICE_X158Y124_A5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_BMUX = CLBLM_R_X101Y124_SLICE_X158Y124_B5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_CMUX = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A = CLBLM_R_X101Y124_SLICE_X159Y124_AO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B = CLBLM_R_X101Y124_SLICE_X159Y124_BO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C = CLBLM_R_X101Y124_SLICE_X159Y124_CO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D = CLBLM_R_X101Y124_SLICE_X159Y124_DO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_AMUX = CLBLM_R_X101Y124_SLICE_X159Y124_A5Q;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A = CLBLM_R_X101Y125_SLICE_X158Y125_AO6;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B = CLBLM_R_X101Y125_SLICE_X158Y125_BO6;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C = CLBLM_R_X101Y125_SLICE_X158Y125_CO6;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D = CLBLM_R_X101Y125_SLICE_X158Y125_DO6;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_BMUX = CLBLM_R_X101Y125_SLICE_X158Y125_B5Q;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A = CLBLM_R_X101Y125_SLICE_X159Y125_AO6;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B = CLBLM_R_X101Y125_SLICE_X159Y125_BO6;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C = CLBLM_R_X101Y125_SLICE_X159Y125_CO6;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D = CLBLM_R_X101Y125_SLICE_X159Y125_DO6;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A = CLBLM_R_X101Y126_SLICE_X158Y126_AO6;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B = CLBLM_R_X101Y126_SLICE_X158Y126_BO6;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C = CLBLM_R_X101Y126_SLICE_X158Y126_CO6;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D = CLBLM_R_X101Y126_SLICE_X158Y126_DO6;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_AMUX = CLBLM_R_X101Y126_SLICE_X158Y126_A5Q;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A = CLBLM_R_X101Y126_SLICE_X159Y126_AO6;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B = CLBLM_R_X101Y126_SLICE_X159Y126_BO6;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C = CLBLM_R_X101Y126_SLICE_X159Y126_CO6;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D = CLBLM_R_X101Y126_SLICE_X159Y126_DO6;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_AMUX = CLBLM_R_X101Y126_SLICE_X159Y126_A5Q;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A = CLBLM_R_X101Y127_SLICE_X158Y127_AO6;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B = CLBLM_R_X101Y127_SLICE_X158Y127_BO6;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C = CLBLM_R_X101Y127_SLICE_X158Y127_CO6;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D = CLBLM_R_X101Y127_SLICE_X158Y127_DO6;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A = CLBLM_R_X101Y127_SLICE_X159Y127_AO6;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B = CLBLM_R_X101Y127_SLICE_X159Y127_BO6;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C = CLBLM_R_X101Y127_SLICE_X159Y127_CO6;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D = CLBLM_R_X101Y127_SLICE_X159Y127_DO6;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_AMUX = CLBLM_R_X101Y127_SLICE_X159Y127_A5Q;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A = CLBLM_R_X101Y128_SLICE_X158Y128_AO6;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B = CLBLM_R_X101Y128_SLICE_X158Y128_BO6;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C = CLBLM_R_X101Y128_SLICE_X158Y128_CO6;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D = CLBLM_R_X101Y128_SLICE_X158Y128_DO6;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_AMUX = CLBLM_R_X101Y128_SLICE_X158Y128_A5Q;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A = CLBLM_R_X101Y128_SLICE_X159Y128_AO6;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B = CLBLM_R_X101Y128_SLICE_X159Y128_BO6;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C = CLBLM_R_X101Y128_SLICE_X159Y128_CO6;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D = CLBLM_R_X101Y128_SLICE_X159Y128_DO6;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A = CLBLM_R_X101Y129_SLICE_X158Y129_AO6;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B = CLBLM_R_X101Y129_SLICE_X158Y129_BO6;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C = CLBLM_R_X101Y129_SLICE_X158Y129_CO6;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D = CLBLM_R_X101Y129_SLICE_X158Y129_DO6;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_AMUX = CLBLM_R_X101Y129_SLICE_X158Y129_A5Q;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_BMUX = CLBLM_R_X101Y129_SLICE_X158Y129_B5Q;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A = CLBLM_R_X101Y129_SLICE_X159Y129_AO6;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B = CLBLM_R_X101Y129_SLICE_X159Y129_BO6;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C = CLBLM_R_X101Y129_SLICE_X159Y129_CO6;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D = CLBLM_R_X101Y129_SLICE_X159Y129_DO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A = CLBLM_R_X101Y130_SLICE_X158Y130_AO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B = CLBLM_R_X101Y130_SLICE_X158Y130_BO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C = CLBLM_R_X101Y130_SLICE_X158Y130_CO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D = CLBLM_R_X101Y130_SLICE_X158Y130_DO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_AMUX = CLBLM_R_X101Y130_SLICE_X158Y130_A5Q;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_CMUX = CLBLM_R_X101Y130_SLICE_X158Y130_C5Q;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A = CLBLM_R_X101Y130_SLICE_X159Y130_AO6;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B = CLBLM_R_X101Y130_SLICE_X159Y130_BO6;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C = CLBLM_R_X101Y130_SLICE_X159Y130_CO6;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D = CLBLM_R_X101Y130_SLICE_X159Y130_DO6;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_BMUX = CLBLM_R_X101Y130_SLICE_X159Y130_B5Q;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_CMUX = CLBLM_R_X101Y130_SLICE_X159Y130_CO6;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A = CLBLM_R_X101Y131_SLICE_X158Y131_AO6;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B = CLBLM_R_X101Y131_SLICE_X158Y131_BO6;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C = CLBLM_R_X101Y131_SLICE_X158Y131_CO6;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D = CLBLM_R_X101Y131_SLICE_X158Y131_DO6;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_BMUX = CLBLM_R_X101Y131_SLICE_X158Y131_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_CMUX = CLBLM_R_X101Y131_SLICE_X158Y131_CO6;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A = CLBLM_R_X101Y131_SLICE_X159Y131_AO6;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B = CLBLM_R_X101Y131_SLICE_X159Y131_BO6;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C = CLBLM_R_X101Y131_SLICE_X159Y131_CO6;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D = CLBLM_R_X101Y131_SLICE_X159Y131_DO6;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_AMUX = CLBLM_R_X101Y131_SLICE_X159Y131_A5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_BMUX = CLBLM_R_X101Y131_SLICE_X159Y131_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_CMUX = CLBLM_R_X101Y131_SLICE_X159Y131_C5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_DMUX = CLBLM_R_X101Y131_SLICE_X159Y131_D5Q;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A = CLBLM_R_X101Y132_SLICE_X158Y132_AO6;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B = CLBLM_R_X101Y132_SLICE_X158Y132_BO6;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C = CLBLM_R_X101Y132_SLICE_X158Y132_CO6;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D = CLBLM_R_X101Y132_SLICE_X158Y132_DO6;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_AMUX = CLBLM_R_X101Y132_SLICE_X158Y132_A5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A = CLBLM_R_X101Y132_SLICE_X159Y132_AO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B = CLBLM_R_X101Y132_SLICE_X159Y132_BO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C = CLBLM_R_X101Y132_SLICE_X159Y132_CO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D = CLBLM_R_X101Y132_SLICE_X159Y132_DO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_BMUX = CLBLM_R_X101Y132_SLICE_X159Y132_B5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_CMUX = CLBLM_R_X101Y132_SLICE_X159Y132_CO6;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A = CLBLM_R_X101Y133_SLICE_X158Y133_AO6;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B = CLBLM_R_X101Y133_SLICE_X158Y133_BO6;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C = CLBLM_R_X101Y133_SLICE_X158Y133_CO6;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D = CLBLM_R_X101Y133_SLICE_X158Y133_DO6;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_BMUX = CLBLM_R_X101Y133_SLICE_X158Y133_B5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A = CLBLM_R_X101Y133_SLICE_X159Y133_AO6;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B = CLBLM_R_X101Y133_SLICE_X159Y133_BO6;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C = CLBLM_R_X101Y133_SLICE_X159Y133_CO6;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D = CLBLM_R_X101Y133_SLICE_X159Y133_DO6;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_AMUX = CLBLM_R_X101Y133_SLICE_X159Y133_A5Q;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A = CLBLM_R_X101Y134_SLICE_X158Y134_AO6;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B = CLBLM_R_X101Y134_SLICE_X158Y134_BO6;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C = CLBLM_R_X101Y134_SLICE_X158Y134_CO6;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D = CLBLM_R_X101Y134_SLICE_X158Y134_DO6;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_AMUX = CLBLM_R_X101Y134_SLICE_X158Y134_A5Q;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A = CLBLM_R_X101Y134_SLICE_X159Y134_AO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B = CLBLM_R_X101Y134_SLICE_X159Y134_BO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C = CLBLM_R_X101Y134_SLICE_X159Y134_CO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D = CLBLM_R_X101Y134_SLICE_X159Y134_DO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_CMUX = CLBLM_R_X101Y134_SLICE_X159Y134_C5Q;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A = CLBLM_R_X101Y135_SLICE_X158Y135_AO6;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B = CLBLM_R_X101Y135_SLICE_X158Y135_BO6;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C = CLBLM_R_X101Y135_SLICE_X158Y135_CO6;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D = CLBLM_R_X101Y135_SLICE_X158Y135_DO6;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_AMUX = CLBLM_R_X101Y135_SLICE_X158Y135_A5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A = CLBLM_R_X101Y135_SLICE_X159Y135_AO6;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B = CLBLM_R_X101Y135_SLICE_X159Y135_BO6;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C = CLBLM_R_X101Y135_SLICE_X159Y135_CO6;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D = CLBLM_R_X101Y135_SLICE_X159Y135_DO6;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_AMUX = CLBLM_R_X101Y135_SLICE_X159Y135_A5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_BMUX = CLBLM_R_X101Y135_SLICE_X159Y135_B5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_CMUX = CLBLM_R_X101Y135_SLICE_X159Y135_C5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_DMUX = CLBLM_R_X101Y135_SLICE_X159Y135_D5Q;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A = CLBLM_R_X101Y136_SLICE_X158Y136_AO6;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B = CLBLM_R_X101Y136_SLICE_X158Y136_BO6;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C = CLBLM_R_X101Y136_SLICE_X158Y136_CO6;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D = CLBLM_R_X101Y136_SLICE_X158Y136_DO6;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_AMUX = CLBLM_R_X101Y136_SLICE_X158Y136_A5Q;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A = CLBLM_R_X101Y136_SLICE_X159Y136_AO6;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B = CLBLM_R_X101Y136_SLICE_X159Y136_BO6;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C = CLBLM_R_X101Y136_SLICE_X159Y136_CO6;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D = CLBLM_R_X101Y136_SLICE_X159Y136_DO6;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_BMUX = CLBLM_R_X101Y136_SLICE_X159Y136_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A = CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B = CLBLM_R_X103Y111_SLICE_X162Y111_BO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C = CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D = CLBLM_R_X103Y111_SLICE_X162Y111_DO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_AMUX = CLBLM_R_X103Y111_SLICE_X162Y111_AO5;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_BMUX = CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_CMUX = CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A = CLBLM_R_X103Y111_SLICE_X163Y111_AO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B = CLBLM_R_X103Y111_SLICE_X163Y111_BO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C = CLBLM_R_X103Y111_SLICE_X163Y111_CO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D = CLBLM_R_X103Y111_SLICE_X163Y111_DO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A = CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B = CLBLM_R_X103Y112_SLICE_X162Y112_BO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C = CLBLM_R_X103Y112_SLICE_X162Y112_CO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D = CLBLM_R_X103Y112_SLICE_X162Y112_DO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_AMUX = CLBLM_R_X103Y112_SLICE_X162Y112_AO5;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_BMUX = CLBLM_R_X103Y112_SLICE_X162Y112_B5Q;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_CMUX = CLBLM_R_X103Y112_SLICE_X162Y112_C5Q;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A = CLBLM_R_X103Y112_SLICE_X163Y112_AO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B = CLBLM_R_X103Y112_SLICE_X163Y112_BO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C = CLBLM_R_X103Y112_SLICE_X163Y112_CO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D = CLBLM_R_X103Y112_SLICE_X163Y112_DO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_AMUX = CLBLM_R_X103Y112_SLICE_X163Y112_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A = CLBLM_R_X103Y113_SLICE_X162Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B = CLBLM_R_X103Y113_SLICE_X162Y113_BO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C = CLBLM_R_X103Y113_SLICE_X162Y113_CO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D = CLBLM_R_X103Y113_SLICE_X162Y113_DO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_AMUX = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_BMUX = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B = CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C = CLBLM_R_X103Y113_SLICE_X163Y113_CO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D = CLBLM_R_X103Y113_SLICE_X163Y113_DO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_BMUX = CLBLM_R_X103Y113_SLICE_X163Y113_BO5;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A = CLBLM_R_X103Y116_SLICE_X162Y116_AO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B = CLBLM_R_X103Y116_SLICE_X162Y116_BO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C = CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_BMUX = CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_DMUX = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A = CLBLM_R_X103Y116_SLICE_X163Y116_AO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B = CLBLM_R_X103Y116_SLICE_X163Y116_BO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D = CLBLM_R_X103Y116_SLICE_X163Y116_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A = CLBLM_R_X103Y117_SLICE_X162Y117_AO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B = CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C = CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D = CLBLM_R_X103Y117_SLICE_X162Y117_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_BMUX = CLBLM_R_X103Y117_SLICE_X162Y117_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A = CLBLM_R_X103Y117_SLICE_X163Y117_AO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B = CLBLM_R_X103Y117_SLICE_X163Y117_BO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C = CLBLM_R_X103Y117_SLICE_X163Y117_CO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D = CLBLM_R_X103Y117_SLICE_X163Y117_DO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A = CLBLM_R_X103Y119_SLICE_X162Y119_AO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B = CLBLM_R_X103Y119_SLICE_X162Y119_BO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C = CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D = CLBLM_R_X103Y119_SLICE_X162Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A = CLBLM_R_X103Y119_SLICE_X163Y119_AO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B = CLBLM_R_X103Y119_SLICE_X163Y119_BO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C = CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D = CLBLM_R_X103Y119_SLICE_X163Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_BMUX = CLBLM_R_X103Y119_SLICE_X163Y119_B5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A = CLBLM_R_X103Y120_SLICE_X162Y120_AO6;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B = CLBLM_R_X103Y120_SLICE_X162Y120_BO6;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C = CLBLM_R_X103Y120_SLICE_X162Y120_CO6;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D = CLBLM_R_X103Y120_SLICE_X162Y120_DO6;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_AMUX = CLBLM_R_X103Y120_SLICE_X162Y120_A5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_BMUX = CLBLM_R_X103Y120_SLICE_X162Y120_B5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_CMUX = CLBLM_R_X103Y120_SLICE_X162Y120_C5Q;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A = CLBLM_R_X103Y120_SLICE_X163Y120_AO6;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B = CLBLM_R_X103Y120_SLICE_X163Y120_BO6;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C = CLBLM_R_X103Y120_SLICE_X163Y120_CO6;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D = CLBLM_R_X103Y120_SLICE_X163Y120_DO6;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_BMUX = CLBLM_R_X103Y120_SLICE_X163Y120_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A = CLBLM_R_X103Y121_SLICE_X162Y121_AO6;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B = CLBLM_R_X103Y121_SLICE_X162Y121_BO6;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C = CLBLM_R_X103Y121_SLICE_X162Y121_CO6;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D = CLBLM_R_X103Y121_SLICE_X162Y121_DO6;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_BMUX = CLBLM_R_X103Y121_SLICE_X162Y121_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A = CLBLM_R_X103Y121_SLICE_X163Y121_AO6;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B = CLBLM_R_X103Y121_SLICE_X163Y121_BO6;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C = CLBLM_R_X103Y121_SLICE_X163Y121_CO6;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D = CLBLM_R_X103Y121_SLICE_X163Y121_DO6;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_AMUX = CLBLM_R_X103Y121_SLICE_X163Y121_A5Q;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_BMUX = CLBLM_R_X103Y121_SLICE_X163Y121_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_CMUX = CLBLM_R_X103Y121_SLICE_X163Y121_C5Q;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A = CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B = CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C = CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D = CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_AMUX = CLBLM_R_X103Y122_SLICE_X162Y122_A5Q;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_BMUX = CLBLM_R_X103Y122_SLICE_X162Y122_B5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_AMUX = CLBLM_R_X103Y122_SLICE_X163Y122_A5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_BMUX = CLBLM_R_X103Y122_SLICE_X163Y122_B5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_CMUX = CLBLM_R_X103Y122_SLICE_X163Y122_C5Q;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A = CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B = CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C = CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D = CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_AMUX = CLBLM_R_X103Y123_SLICE_X162Y123_A5Q;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A = CLBLM_R_X103Y123_SLICE_X163Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B = CLBLM_R_X103Y123_SLICE_X163Y123_BO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C = CLBLM_R_X103Y123_SLICE_X163Y123_CO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D = CLBLM_R_X103Y123_SLICE_X163Y123_DO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A = CLBLM_R_X103Y124_SLICE_X162Y124_AO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B = CLBLM_R_X103Y124_SLICE_X162Y124_BO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C = CLBLM_R_X103Y124_SLICE_X162Y124_CO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D = CLBLM_R_X103Y124_SLICE_X162Y124_DO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_BMUX = CLBLM_R_X103Y124_SLICE_X162Y124_B5Q;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_DMUX = CLBLM_R_X103Y124_SLICE_X162Y124_DO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A = CLBLM_R_X103Y124_SLICE_X163Y124_AO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B = CLBLM_R_X103Y124_SLICE_X163Y124_BO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C = CLBLM_R_X103Y124_SLICE_X163Y124_CO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D = CLBLM_R_X103Y124_SLICE_X163Y124_DO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_BMUX = CLBLM_R_X103Y124_SLICE_X163Y124_B5Q;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_DMUX = CLBLM_R_X103Y124_SLICE_X163Y124_DO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A = CLBLM_R_X103Y125_SLICE_X162Y125_AO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B = CLBLM_R_X103Y125_SLICE_X162Y125_BO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C = CLBLM_R_X103Y125_SLICE_X162Y125_CO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D = CLBLM_R_X103Y125_SLICE_X162Y125_DO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_AMUX = CLBLM_R_X103Y125_SLICE_X162Y125_A5Q;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_CMUX = CLBLM_R_X103Y125_SLICE_X162Y125_C5Q;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A = CLBLM_R_X103Y125_SLICE_X163Y125_AO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B = CLBLM_R_X103Y125_SLICE_X163Y125_BO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C = CLBLM_R_X103Y125_SLICE_X163Y125_CO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D = CLBLM_R_X103Y125_SLICE_X163Y125_DO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_BMUX = CLBLM_R_X103Y125_SLICE_X163Y125_B5Q;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_CMUX = CLBLM_R_X103Y125_SLICE_X163Y125_C5Q;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A = CLBLM_R_X103Y126_SLICE_X162Y126_AO6;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B = CLBLM_R_X103Y126_SLICE_X162Y126_BO6;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C = CLBLM_R_X103Y126_SLICE_X162Y126_CO6;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D = CLBLM_R_X103Y126_SLICE_X162Y126_DO6;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_BMUX = CLBLM_R_X103Y126_SLICE_X162Y126_B5Q;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A = CLBLM_R_X103Y126_SLICE_X163Y126_AO6;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B = CLBLM_R_X103Y126_SLICE_X163Y126_BO6;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C = CLBLM_R_X103Y126_SLICE_X163Y126_CO6;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D = CLBLM_R_X103Y126_SLICE_X163Y126_DO6;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_AMUX = CLBLM_R_X103Y126_SLICE_X163Y126_A5Q;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A = CLBLM_R_X103Y127_SLICE_X162Y127_AO6;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B = CLBLM_R_X103Y127_SLICE_X162Y127_BO6;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C = CLBLM_R_X103Y127_SLICE_X162Y127_CO6;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D = CLBLM_R_X103Y127_SLICE_X162Y127_DO6;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A = CLBLM_R_X103Y127_SLICE_X163Y127_AO6;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B = CLBLM_R_X103Y127_SLICE_X163Y127_BO6;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C = CLBLM_R_X103Y127_SLICE_X163Y127_CO6;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D = CLBLM_R_X103Y127_SLICE_X163Y127_DO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_OQ = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y5_OLOGIC_X0Y6_OQ = 1'b0;
  assign LIOI3_X0Y5_OLOGIC_X0Y6_TQ = 1'b1;
  assign LIOI3_X0Y5_OLOGIC_X0Y5_OQ = 1'b0;
  assign LIOI3_X0Y5_OLOGIC_X0Y5_TQ = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_OQ = 1'b0;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_TQ = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_OQ = 1'b0;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_TQ = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_OQ = 1'b0;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_TQ = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_OQ = 1'b0;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_TQ = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_OQ = 1'b0;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_TQ = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_OQ = 1'b0;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_OQ = 1'b0;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_OQ = 1'b0;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_TQ = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_OQ = 1'b0;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_TQ = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_OQ = 1'b0;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = 1'b0;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = 1'b0;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_OQ = 1'b0;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_TQ = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_OQ = 1'b0;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_TQ = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_OQ = 1'b0;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_TQ = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_OQ = 1'b0;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_TQ = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_OQ = 1'b0;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_TQ = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_OQ = 1'b0;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_TQ = 1'b1;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_OQ = 1'b0;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_TQ = 1'b1;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_OQ = 1'b0;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_TQ = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_OQ = 1'b0;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_TQ = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_OQ = 1'b0;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_TQ = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = 1'b0;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_OQ = 1'b0;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_TQ = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_OQ = 1'b0;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_TQ = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_OQ = 1'b0;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_TQ = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_OQ = 1'b0;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_TQ = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_OQ = 1'b0;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_TQ = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_OQ = 1'b0;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_TQ = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_OQ = 1'b0;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_TQ = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_OQ = 1'b0;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_TQ = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_OQ = 1'b0;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_TQ = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_OQ = 1'b0;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_TQ = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_OQ = 1'b0;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_TQ = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_OQ = 1'b0;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_TQ = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_OQ = 1'b0;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = 1'b0;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = 1'b0;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = 1'b0;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = 1'b0;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = 1'b0;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = 1'b0;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = 1'b0;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = 1'b0;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = 1'b0;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = 1'b0;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = 1'b0;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = 1'b0;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = 1'b0;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = 1'b0;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = 1'b0;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = 1'b0;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = 1'b0;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = 1'b0;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = 1'b0;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = 1'b0;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = 1'b0;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = 1'b0;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = 1'b0;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = 1'b0;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = 1'b0;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = 1'b0;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = 1'b0;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = 1'b0;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = 1'b0;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = 1'b0;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = 1'b0;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = 1'b0;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = 1'b0;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = 1'b0;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = 1'b0;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = 1'b0;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = 1'b0;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = 1'b0;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = 1'b0;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = 1'b0;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = 1'b0;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = 1'b0;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = 1'b0;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = 1'b0;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = 1'b0;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = 1'b0;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = 1'b0;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = 1'b0;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = 1'b0;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = 1'b0;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = 1'b0;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = 1'b0;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = 1'b0;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = 1'b0;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = 1'b0;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = 1'b0;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b0;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = 1'b0;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_X0Y201_OLOGIC_X0Y202_OQ = 1'b0;
  assign LIOI3_X0Y201_OLOGIC_X0Y202_TQ = 1'b1;
  assign LIOI3_X0Y201_OLOGIC_X0Y201_OQ = 1'b0;
  assign LIOI3_X0Y201_OLOGIC_X0Y201_TQ = 1'b1;
  assign LIOI3_X0Y203_OLOGIC_X0Y204_OQ = 1'b0;
  assign LIOI3_X0Y203_OLOGIC_X0Y204_TQ = 1'b1;
  assign LIOI3_X0Y203_OLOGIC_X0Y203_OQ = 1'b0;
  assign LIOI3_X0Y203_OLOGIC_X0Y203_TQ = 1'b1;
  assign LIOI3_X0Y205_OLOGIC_X0Y206_OQ = 1'b0;
  assign LIOI3_X0Y205_OLOGIC_X0Y206_TQ = 1'b1;
  assign LIOI3_X0Y205_OLOGIC_X0Y205_OQ = 1'b0;
  assign LIOI3_X0Y205_OLOGIC_X0Y205_TQ = 1'b1;
  assign LIOI3_X0Y209_OLOGIC_X0Y210_OQ = 1'b0;
  assign LIOI3_X0Y209_OLOGIC_X0Y210_TQ = 1'b1;
  assign LIOI3_X0Y209_OLOGIC_X0Y209_OQ = 1'b0;
  assign LIOI3_X0Y209_OLOGIC_X0Y209_TQ = 1'b1;
  assign LIOI3_X0Y211_OLOGIC_X0Y212_OQ = 1'b0;
  assign LIOI3_X0Y211_OLOGIC_X0Y212_TQ = 1'b1;
  assign LIOI3_X0Y211_OLOGIC_X0Y211_OQ = 1'b0;
  assign LIOI3_X0Y211_OLOGIC_X0Y211_TQ = 1'b1;
  assign LIOI3_X0Y215_OLOGIC_X0Y216_OQ = 1'b0;
  assign LIOI3_X0Y215_OLOGIC_X0Y216_TQ = 1'b1;
  assign LIOI3_X0Y215_OLOGIC_X0Y215_OQ = 1'b0;
  assign LIOI3_X0Y215_OLOGIC_X0Y215_TQ = 1'b1;
  assign LIOI3_X0Y217_OLOGIC_X0Y218_OQ = 1'b0;
  assign LIOI3_X0Y217_OLOGIC_X0Y218_TQ = 1'b1;
  assign LIOI3_X0Y217_OLOGIC_X0Y217_OQ = 1'b0;
  assign LIOI3_X0Y217_OLOGIC_X0Y217_TQ = 1'b1;
  assign LIOI3_X0Y221_OLOGIC_X0Y222_OQ = 1'b0;
  assign LIOI3_X0Y221_OLOGIC_X0Y222_TQ = 1'b1;
  assign LIOI3_X0Y221_OLOGIC_X0Y221_OQ = 1'b0;
  assign LIOI3_X0Y221_OLOGIC_X0Y221_TQ = 1'b1;
  assign LIOI3_X0Y223_OLOGIC_X0Y224_OQ = 1'b0;
  assign LIOI3_X0Y223_OLOGIC_X0Y224_TQ = 1'b1;
  assign LIOI3_X0Y223_OLOGIC_X0Y223_OQ = 1'b0;
  assign LIOI3_X0Y223_OLOGIC_X0Y223_TQ = 1'b1;
  assign LIOI3_X0Y225_OLOGIC_X0Y226_OQ = 1'b0;
  assign LIOI3_X0Y225_OLOGIC_X0Y226_TQ = 1'b1;
  assign LIOI3_X0Y225_OLOGIC_X0Y225_OQ = 1'b0;
  assign LIOI3_X0Y225_OLOGIC_X0Y225_TQ = 1'b1;
  assign LIOI3_X0Y227_OLOGIC_X0Y228_OQ = 1'b0;
  assign LIOI3_X0Y227_OLOGIC_X0Y228_TQ = 1'b1;
  assign LIOI3_X0Y227_OLOGIC_X0Y227_OQ = 1'b0;
  assign LIOI3_X0Y227_OLOGIC_X0Y227_TQ = 1'b1;
  assign LIOI3_X0Y229_OLOGIC_X0Y230_OQ = 1'b0;
  assign LIOI3_X0Y229_OLOGIC_X0Y230_TQ = 1'b1;
  assign LIOI3_X0Y229_OLOGIC_X0Y229_OQ = 1'b0;
  assign LIOI3_X0Y229_OLOGIC_X0Y229_TQ = 1'b1;
  assign LIOI3_X0Y233_OLOGIC_X0Y234_OQ = 1'b0;
  assign LIOI3_X0Y233_OLOGIC_X0Y234_TQ = 1'b1;
  assign LIOI3_X0Y233_OLOGIC_X0Y233_OQ = 1'b0;
  assign LIOI3_X0Y233_OLOGIC_X0Y233_TQ = 1'b1;
  assign LIOI3_X0Y235_OLOGIC_X0Y236_OQ = 1'b0;
  assign LIOI3_X0Y235_OLOGIC_X0Y236_TQ = 1'b1;
  assign LIOI3_X0Y235_OLOGIC_X0Y235_OQ = 1'b0;
  assign LIOI3_X0Y235_OLOGIC_X0Y235_TQ = 1'b1;
  assign LIOI3_X0Y239_OLOGIC_X0Y240_OQ = 1'b0;
  assign LIOI3_X0Y239_OLOGIC_X0Y240_TQ = 1'b1;
  assign LIOI3_X0Y239_OLOGIC_X0Y239_OQ = 1'b0;
  assign LIOI3_X0Y239_OLOGIC_X0Y239_TQ = 1'b1;
  assign LIOI3_X0Y241_OLOGIC_X0Y242_OQ = 1'b0;
  assign LIOI3_X0Y241_OLOGIC_X0Y242_TQ = 1'b1;
  assign LIOI3_X0Y241_OLOGIC_X0Y241_OQ = 1'b0;
  assign LIOI3_X0Y241_OLOGIC_X0Y241_TQ = 1'b1;
  assign LIOI3_X0Y245_OLOGIC_X0Y246_OQ = 1'b0;
  assign LIOI3_X0Y245_OLOGIC_X0Y246_TQ = 1'b1;
  assign LIOI3_X0Y245_OLOGIC_X0Y245_OQ = 1'b0;
  assign LIOI3_X0Y245_OLOGIC_X0Y245_TQ = 1'b1;
  assign LIOI3_X0Y247_OLOGIC_X0Y248_OQ = 1'b0;
  assign LIOI3_X0Y247_OLOGIC_X0Y248_TQ = 1'b1;
  assign LIOI3_X0Y247_OLOGIC_X0Y247_OQ = 1'b0;
  assign LIOI3_X0Y247_OLOGIC_X0Y247_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ = 1'b0;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_OQ = 1'b0;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_TQ = 1'b1;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_OQ = 1'b0;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = 1'b0;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = 1'b0;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = 1'b0;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b0;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_OQ = 1'b0;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_TQ = 1'b1;
  assign LIOI3_SING_X0Y249_OLOGIC_X0Y249_OQ = 1'b0;
  assign LIOI3_SING_X0Y249_OLOGIC_X0Y249_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_OQ = 1'b0;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_OQ = 1'b0;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_OQ = 1'b0;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_OQ = 1'b0;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_OQ = 1'b0;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_OQ = 1'b0;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_OQ = 1'b0;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_OQ = 1'b0;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_OQ = 1'b0;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_OQ = 1'b0;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_OQ = 1'b0;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_OQ = 1'b0;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_OQ = 1'b0;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_OQ = 1'b0;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_OQ = 1'b0;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_OQ = 1'b0;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_OQ = 1'b0;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_OQ = 1'b0;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_OQ = 1'b0;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_OQ = 1'b0;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_X105Y77_ILOGIC_X1Y78_O = RIOB33_X105Y77_IOB_X1Y78_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_OQ = 1'b0;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_OQ = CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_OQ = 1'b0;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_OQ = CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_OQ = CLBLL_L_X102Y117_SLICE_X160Y117_CO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_OQ = CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_OQ = CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_OQ = CLBLL_L_X102Y116_SLICE_X160Y116_AO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_OQ = CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_OQ = CLBLL_L_X102Y119_SLICE_X160Y119_CO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_OQ = CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_OQ = CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_OQ = CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_OQ = CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_OQ = CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_OQ = 1'b0;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_OQ = 1'b0;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_OQ = 1'b0;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_OQ = 1'b0;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_OQ = 1'b0;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_OQ = 1'b0;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = CLBLM_R_X101Y113_SLICE_X159Y113_AO6;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLM_R_X103Y121_SLICE_X162Y121_CO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = CLBLM_R_X101Y113_SLICE_X159Y113_BO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b0;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b0;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b0;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b0;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = 1'b0;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b0;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = 1'b0;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = 1'b0;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = 1'b0;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = 1'b0;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = 1'b0;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = 1'b0;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = 1'b0;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = 1'b0;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = 1'b0;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = 1'b0;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = 1'b0;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = 1'b0;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = 1'b0;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = 1'b0;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = 1'b0;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = 1'b0;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = 1'b0;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = 1'b0;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = 1'b0;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = 1'b0;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_R_X103Y124_SLICE_X162Y124_CO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLL_L_X102Y120_SLICE_X161Y120_CO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X103Y124_SLICE_X163Y124_CO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLL_L_X102Y124_SLICE_X161Y124_CO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ = 1'b0;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ = CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ = 1'b0;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b0;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLL_L_X102Y123_SLICE_X160Y123_CO6;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ = CLBLM_R_X101Y120_SLICE_X159Y120_CO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ = CLBLL_L_X102Y119_SLICE_X161Y119_CO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ = CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X103Y120_SLICE_X163Y120_CO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLL_L_X102Y118_SLICE_X160Y118_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ = CLBLM_R_X101Y117_SLICE_X159Y117_AO5;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ = CLBLL_L_X100Y115_SLICE_X157Y115_CO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_T1 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = 1'b0;
  assign LIOB33_X0Y147_IOB_X0Y147_O = 1'b0;
  assign LIOB33_X0Y147_IOB_X0Y148_T = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_T = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A2 = CLBLM_R_X97Y112_SLICE_X153Y112_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A3 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A4 = CLBLM_L_X98Y115_SLICE_X154Y115_AQ;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A5 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_A6 = 1'b1;
  assign LIOI3_X0Y217_OLOGIC_X0Y218_D1 = 1'b0;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B2 = CLBLM_R_X95Y111_SLICE_X151Y111_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B3 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B4 = CLBLM_R_X97Y115_SLICE_X153Y115_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B5 = CLBLM_R_X97Y112_SLICE_X153Y112_CO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_B6 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C1 = CLBLL_L_X100Y111_SLICE_X157Y111_C5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C2 = CLBLM_R_X95Y111_SLICE_X151Y111_CO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C4 = CLBLM_R_X97Y112_SLICE_X153Y112_A5Q;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C5 = CLBLM_L_X98Y110_SLICE_X154Y110_BO6;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y217_OLOGIC_X0Y218_T1 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y217_OLOGIC_X0Y217_D1 = 1'b0;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D1 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D2 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D3 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D4 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D5 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_D6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_D1 = 1'b0;
  assign CLBLM_R_X97Y112_SLICE_X153Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y217_OLOGIC_X0Y217_T1 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A2 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A3 = CLBLM_R_X97Y112_SLICE_X153Y112_B5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A4 = CLBLM_R_X95Y111_SLICE_X151Y111_B5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A5 = CLBLM_R_X97Y111_SLICE_X153Y111_BO6;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_A6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_T1 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B2 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B3 = CLBLM_R_X95Y112_SLICE_X150Y112_AQ;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B4 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B5 = CLBLM_R_X97Y112_SLICE_X152Y112_C5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_B6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_D1 = 1'b0;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C1 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C2 = CLBLM_R_X97Y112_SLICE_X152Y112_CQ;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C3 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C5 = CLBLM_R_X95Y112_SLICE_X150Y112_BQ;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_C6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_T1 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D1 = CLBLM_R_X97Y112_SLICE_X152Y112_C5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D2 = CLBLM_R_X97Y112_SLICE_X152Y112_CQ;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D3 = 1'b1;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D5 = CLBLM_R_X97Y112_SLICE_X152Y112_B5Q;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_D6 = CLBLM_R_X95Y112_SLICE_X150Y112_BQ;
  assign CLBLM_R_X97Y112_SLICE_X152Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b0;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_T = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A2 = CLBLM_R_X93Y116_SLICE_X146Y116_CO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B3 = CLBLM_L_X94Y127_SLICE_X149Y127_CO6;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = 1'b0;
  assign LIOB33_X0Y151_IOB_X0Y151_O = 1'b0;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLL_L_X102Y123_SLICE_X160Y123_CO6;
  assign LIOB33_X0Y151_IOB_X0Y152_T = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y151_T = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A1 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A2 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A3 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A5 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_A6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B1 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B2 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B3 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B5 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_B6 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C1 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C2 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B3 = CLBLM_L_X92Y129_SLICE_X145Y129_A5Q;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C3 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C5 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_C6 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B4 = CLBLM_L_X92Y129_SLICE_X145Y129_CQ;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B5 = CLBLM_L_X92Y129_SLICE_X145Y129_C5Q;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D1 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D2 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D3 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D5 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X153Y113_D6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A2 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A3 = CLBLM_R_X97Y113_SLICE_X152Y113_AQ;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A5 = CLBLM_R_X97Y112_SLICE_X152Y112_BQ;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_A6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B2 = CLBLM_R_X97Y112_SLICE_X152Y112_BQ;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B3 = CLBLM_R_X97Y113_SLICE_X152Y113_AQ;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B5 = CLBLM_R_X95Y112_SLICE_X150Y112_AQ;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_B6 = CLBLM_R_X97Y113_SLICE_X152Y113_A5Q;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C1 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C2 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C3 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C5 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_C6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D1 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D2 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D3 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D4 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D5 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_D6 = 1'b1;
  assign CLBLM_R_X97Y113_SLICE_X152Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y153_IOB_X0Y154_O = 1'b0;
  assign LIOB33_X0Y153_IOB_X0Y153_O = 1'b0;
  assign LIOB33_X0Y153_IOB_X0Y154_T = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y153_T = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C4 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C5 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A2 = CLBLM_L_X90Y130_SLICE_X142Y130_AQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A4 = CLBLM_L_X90Y131_SLICE_X142Y131_BO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLL_L_X102Y120_SLICE_X161Y120_CO6;
  assign LIOI3_X0Y221_OLOGIC_X0Y222_D1 = 1'b0;
  assign LIOI3_X0Y221_OLOGIC_X0Y222_T1 = 1'b1;
  assign LIOI3_X0Y221_OLOGIC_X0Y221_D1 = 1'b0;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_D1 = 1'b0;
  assign LIOI3_X0Y221_OLOGIC_X0Y221_T1 = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = 1'b0;
  assign LIOB33_X0Y155_IOB_X0Y155_O = 1'b0;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_D1 = 1'b0;
  assign LIOB33_X0Y155_IOB_X0Y156_T = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y155_T = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_T1 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A2 = CLBLM_R_X97Y116_SLICE_X152Y116_A5Q;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A3 = CLBLM_R_X95Y115_SLICE_X150Y115_C5Q;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A4 = CLBLM_L_X98Y113_SLICE_X154Y113_CO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A5 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_A6 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B2 = CLBLM_R_X97Y115_SLICE_X153Y115_BQ;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B3 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B4 = CLBLM_R_X97Y116_SLICE_X153Y116_BQ;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B5 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_B6 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C1 = CLBLM_R_X97Y116_SLICE_X153Y116_DO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C2 = CLBLM_L_X98Y115_SLICE_X155Y115_CQ;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C5 = CLBLM_R_X97Y115_SLICE_X153Y115_DO6;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_C6 = CLBLL_L_X100Y115_SLICE_X156Y115_C5Q;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D2 = CLBLM_R_X97Y116_SLICE_X153Y116_AQ;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D3 = CLBLM_R_X97Y115_SLICE_X153Y115_BQ;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D4 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D5 = CLBLM_R_X97Y115_SLICE_X153Y115_B5Q;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_D6 = CLBLM_R_X97Y116_SLICE_X153Y116_BQ;
  assign CLBLM_R_X97Y115_SLICE_X153Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A2 = CLBLM_L_X94Y115_SLICE_X148Y115_A5Q;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A3 = CLBLM_L_X98Y116_SLICE_X154Y116_AO6;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A4 = CLBLM_L_X98Y114_SLICE_X154Y114_A5Q;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A5 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_A6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B1 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B2 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B3 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B4 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B5 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_B6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C1 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C2 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C3 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C4 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C5 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_C6 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D1 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D2 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D3 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D4 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D5 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_D6 = 1'b1;
  assign CLBLM_R_X97Y115_SLICE_X152Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y157_IOB_X0Y158_O = 1'b0;
  assign LIOB33_X0Y157_IOB_X0Y157_O = 1'b0;
  assign LIOB33_X0Y157_IOB_X0Y158_T = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y157_T = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A2 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A3 = CLBLM_R_X97Y116_SLICE_X152Y116_CO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A4 = CLBLM_R_X97Y115_SLICE_X153Y115_CO6;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A5 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_A6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B2 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B3 = CLBLM_L_X98Y116_SLICE_X155Y116_B5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B4 = CLBLM_R_X97Y116_SLICE_X153Y116_AQ;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B5 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_B6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C1 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C2 = CLBLM_R_X97Y116_SLICE_X153Y116_CQ;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C4 = CLBLM_R_X97Y116_SLICE_X153Y116_A5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C5 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_C6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D1 = CLBLM_R_X97Y116_SLICE_X153Y116_C5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D2 = CLBLM_R_X97Y116_SLICE_X153Y116_CQ;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D3 = CLBLM_R_X97Y116_SLICE_X152Y116_B5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D4 = CLBLM_R_X97Y116_SLICE_X153Y116_A5Q;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_D6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X153Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A1 = CLBLM_R_X97Y116_SLICE_X152Y116_B5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A2 = CLBLM_L_X90Y116_SLICE_X143Y116_C5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A3 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A4 = CLBLM_L_X98Y115_SLICE_X154Y115_CO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_A6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B2 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B3 = CLBLM_R_X97Y116_SLICE_X153Y116_C5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B4 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B5 = CLBLM_R_X95Y115_SLICE_X150Y115_BQ;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_B6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C1 = CLBLM_R_X93Y120_SLICE_X147Y120_DO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C2 = CLBLM_R_X95Y116_SLICE_X151Y116_A5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C3 = CLBLM_R_X97Y116_SLICE_X153Y116_DO6;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C4 = CLBLM_R_X97Y116_SLICE_X152Y116_A5Q;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D1 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D2 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D3 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D4 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D5 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_D6 = 1'b1;
  assign CLBLM_R_X97Y116_SLICE_X152Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = 1'b0;
  assign LIOB33_X0Y159_IOB_X0Y159_O = 1'b0;
  assign LIOB33_X0Y159_IOB_X0Y160_T = 1'b1;
  assign LIOB33_X0Y159_IOB_X0Y159_T = 1'b1;
  assign LIOI3_X0Y223_OLOGIC_X0Y224_D1 = 1'b0;
  assign LIOI3_X0Y223_OLOGIC_X0Y224_T1 = 1'b1;
  assign LIOI3_X0Y223_OLOGIC_X0Y223_D1 = 1'b0;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = 1'b0;
  assign LIOI3_X0Y223_OLOGIC_X0Y223_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = 1'b0;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = 1'b0;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A2 = CLBLM_R_X97Y117_SLICE_X153Y117_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A3 = CLBLM_R_X97Y119_SLICE_X153Y119_AQ;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A4 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A5 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_D1 = 1'b0;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B4 = CLBLM_R_X97Y117_SLICE_X153Y117_DO5;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B5 = CLBLM_L_X90Y116_SLICE_X142Y116_DO6;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_B6 = CLBLM_R_X97Y117_SLICE_X153Y117_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C1 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C2 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C4 = CLBLM_R_X93Y117_SLICE_X146Y117_AQ;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C5 = CLBLM_R_X97Y118_SLICE_X153Y118_BQ;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_T1 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D1 = CLBLM_R_X97Y117_SLICE_X153Y117_C5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D2 = CLBLM_R_X97Y117_SLICE_X153Y117_BQ;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D4 = CLBLM_R_X97Y117_SLICE_X152Y117_B5Q;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D5 = CLBLM_R_X97Y118_SLICE_X153Y118_BQ;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_D6 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X153Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A2 = CLBLM_R_X97Y117_SLICE_X153Y117_CQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A3 = CLBLM_R_X97Y117_SLICE_X152Y117_AQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A4 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A5 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_A6 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B2 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B3 = CLBLL_L_X100Y118_SLICE_X157Y118_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B4 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B5 = CLBLM_R_X95Y117_SLICE_X150Y117_C5Q;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_B6 = CLBLM_R_X97Y117_SLICE_X152Y117_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_BX = CLBLM_R_X97Y117_SLICE_X153Y117_DO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C1 = CLBLM_R_X97Y117_SLICE_X153Y117_AQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C2 = CLBLM_R_X97Y117_SLICE_X152Y117_BQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C3 = CLBLM_R_X89Y115_SLICE_X141Y115_DO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C5 = CLBLM_R_X97Y117_SLICE_X152Y117_DO6;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y161_IOB_X0Y162_O = 1'b0;
  assign LIOB33_X0Y161_IOB_X0Y161_O = 1'b0;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D1 = CLBLM_R_X97Y117_SLICE_X153Y117_CQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D2 = CLBLM_R_X93Y117_SLICE_X146Y117_AQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D3 = CLBLM_R_X97Y117_SLICE_X152Y117_AQ;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D4 = CLBLM_R_X97Y117_SLICE_X152Y117_A5Q;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D5 = 1'b1;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y117_SLICE_X152Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y161_IOB_X0Y161_T = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y162_T = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = 1'b0;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A1 = CLBLM_R_X97Y118_SLICE_X153Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A2 = CLBLM_R_X97Y119_SLICE_X153Y119_BQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A3 = CLBLM_R_X97Y118_SLICE_X153Y118_AQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A4 = CLBLM_R_X97Y118_SLICE_X152Y118_C5Q;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_A6 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B2 = CLBLM_R_X97Y118_SLICE_X152Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B3 = CLBLM_R_X97Y117_SLICE_X153Y117_BQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B4 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B5 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_B6 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C1 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C2 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C4 = CLBLM_R_X97Y119_SLICE_X153Y119_BQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C5 = CLBLM_L_X98Y120_SLICE_X154Y120_CQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_C6 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D2 = CLBLM_R_X97Y118_SLICE_X153Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D3 = CLBLM_R_X97Y119_SLICE_X153Y119_BQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D4 = CLBLL_L_X100Y118_SLICE_X157Y118_B5Q;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D5 = CLBLM_R_X97Y118_SLICE_X153Y118_AQ;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_D6 = CLBLM_R_X97Y118_SLICE_X152Y118_C5Q;
  assign CLBLM_R_X97Y118_SLICE_X153Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A3 = CLBLM_L_X90Y117_SLICE_X142Y117_DO6;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A4 = CLBLM_R_X97Y118_SLICE_X152Y118_BO6;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A5 = CLBLM_R_X97Y119_SLICE_X153Y119_AQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y163_IOB_X0Y163_O = 1'b0;
  assign LIOB33_X0Y163_IOB_X0Y164_O = 1'b0;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_AX = CLBLM_R_X97Y118_SLICE_X152Y118_BO5;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B2 = CLBLM_R_X97Y118_SLICE_X153Y118_B5Q;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B3 = CLBLM_R_X97Y118_SLICE_X152Y118_AQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B4 = CLBLM_R_X97Y118_SLICE_X152Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B5 = CLBLM_R_X97Y118_SLICE_X152Y118_A5Q;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_B6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_T = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y164_T = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C1 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C2 = CLBLM_R_X97Y118_SLICE_X152Y118_AQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C4 = CLBLM_R_X97Y118_SLICE_X153Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C5 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_C6 = 1'b1;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D1 = CLBLM_R_X97Y118_SLICE_X152Y118_A5Q;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D2 = CLBLM_R_X97Y118_SLICE_X152Y118_AQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D3 = CLBLM_R_X97Y118_SLICE_X153Y118_B5Q;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D4 = CLBLL_L_X100Y118_SLICE_X157Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_D6 = CLBLM_R_X97Y118_SLICE_X152Y118_CQ;
  assign CLBLM_R_X97Y118_SLICE_X152Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C1 = CLBLM_L_X90Y126_SLICE_X142Y126_CQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOB33_X0Y55_IOB_X0Y56_T = 1'b1;
  assign LIOB33_X0Y55_IOB_X0Y55_T = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A2 = CLBLM_R_X97Y119_SLICE_X153Y119_A5Q;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A3 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A4 = CLBLM_L_X98Y119_SLICE_X154Y119_AQ;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A5 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_A6 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B2 = CLBLM_R_X97Y119_SLICE_X153Y119_A5Q;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B5 = CLBLM_R_X97Y118_SLICE_X153Y118_AO6;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_B6 = CLBLM_L_X90Y119_SLICE_X142Y119_DO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = 1'b0;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C1 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C2 = CLBLM_R_X97Y119_SLICE_X153Y119_CQ;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C4 = CLBLM_R_X97Y120_SLICE_X153Y120_BQ;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C5 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_C6 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y165_O = 1'b0;
  assign LIOB33_X0Y165_IOB_X0Y166_O = 1'b0;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y165_IOB_X0Y165_T = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D1 = CLBLM_R_X97Y119_SLICE_X153Y119_C5Q;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D2 = CLBLM_R_X97Y119_SLICE_X153Y119_CQ;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D4 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D5 = CLBLM_R_X95Y119_SLICE_X150Y119_B5Q;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_D6 = CLBLM_R_X97Y120_SLICE_X153Y120_BQ;
  assign LIOB33_X0Y165_IOB_X0Y166_T = 1'b1;
  assign LIOI3_X0Y225_OLOGIC_X0Y226_D1 = 1'b0;
  assign CLBLM_R_X97Y119_SLICE_X153Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y225_OLOGIC_X0Y226_T1 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A2 = CLBLM_R_X97Y119_SLICE_X152Y119_A5Q;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A3 = CLBLL_L_X100Y122_SLICE_X156Y122_AQ;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A4 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A5 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_A6 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B1 = CLBLM_R_X97Y119_SLICE_X152Y119_DO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B3 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B4 = CLBLM_L_X98Y120_SLICE_X154Y120_DO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B5 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_B6 = 1'b1;
  assign LIOI3_X0Y225_OLOGIC_X0Y225_D1 = 1'b0;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = 1'b0;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C1 = CLBLL_L_X100Y119_SLICE_X156Y119_AQ;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C2 = CLBLL_L_X100Y118_SLICE_X157Y118_A5Q;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C4 = CLBLM_R_X97Y120_SLICE_X152Y120_BQ;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C5 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_C6 = 1'b1;
  assign LIOI3_X0Y225_OLOGIC_X0Y225_T1 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D2 = CLBLM_R_X95Y118_SLICE_X151Y118_CO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D3 = CLBLM_R_X97Y119_SLICE_X152Y119_AQ;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D4 = CLBLM_L_X98Y119_SLICE_X155Y119_DO6;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_D6 = CLBLM_R_X95Y118_SLICE_X150Y118_A5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = 1'b0;
  assign CLBLM_R_X97Y119_SLICE_X152Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_D1 = 1'b0;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_D1 = 1'b0;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_T1 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = 1'b0;
  assign LIOB33_X0Y167_IOB_X0Y167_O = 1'b0;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A1 = CLBLM_R_X97Y120_SLICE_X153Y120_B5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A3 = CLBLM_L_X98Y120_SLICE_X155Y120_B5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A4 = CLBLM_R_X97Y120_SLICE_X152Y120_CO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A5 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_A6 = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y167_T = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y168_T = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B2 = CLBLM_L_X98Y120_SLICE_X155Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B3 = CLBLL_L_X102Y121_SLICE_X161Y121_C5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B4 = CLBLM_R_X97Y120_SLICE_X152Y120_DO6;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B5 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_B6 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C1 = CLBLL_L_X100Y120_SLICE_X157Y120_BQ;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C2 = CLBLL_L_X100Y118_SLICE_X157Y118_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C4 = CLBLM_R_X97Y121_SLICE_X153Y121_CQ;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C5 = CLBLL_L_X100Y119_SLICE_X157Y119_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_C6 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D1 = CLBLL_L_X102Y121_SLICE_X160Y121_AQ;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D2 = CLBLM_R_X97Y120_SLICE_X153Y120_CQ;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D3 = CLBLM_R_X97Y120_SLICE_X153Y120_DQ;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D4 = CLBLM_R_X101Y120_SLICE_X158Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_D6 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X153Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A2 = CLBLM_R_X97Y120_SLICE_X152Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A3 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A4 = CLBLM_R_X97Y119_SLICE_X152Y119_AQ;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A5 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_A6 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B2 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B3 = CLBLM_R_X97Y123_SLICE_X152Y123_C5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B4 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B5 = 1'b1;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_B6 = CLBLM_L_X98Y120_SLICE_X154Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C1 = CLBLM_L_X94Y119_SLICE_X149Y119_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C2 = CLBLM_R_X97Y120_SLICE_X152Y120_AQ;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C4 = CLBLM_L_X98Y124_SLICE_X154Y124_DO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_C6 = CLBLM_R_X95Y119_SLICE_X150Y119_DO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D1 = CLBLM_L_X98Y120_SLICE_X155Y120_DO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D3 = CLBLM_R_X97Y119_SLICE_X153Y119_DO6;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D4 = CLBLM_R_X97Y120_SLICE_X152Y120_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_D6 = CLBLM_R_X95Y119_SLICE_X150Y119_A5Q;
  assign CLBLM_R_X97Y120_SLICE_X152Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y169_IOB_X0Y170_O = 1'b0;
  assign LIOB33_X0Y169_IOB_X0Y169_O = 1'b0;
  assign LIOB33_X0Y169_IOB_X0Y170_T = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_T = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A2 = CLBLM_R_X97Y120_SLICE_X152Y120_AQ;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A3 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A4 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A5 = CLBLM_R_X97Y121_SLICE_X153Y121_A5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_A6 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B2 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B3 = CLBLM_L_X98Y124_SLICE_X154Y124_A5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B4 = CLBLM_R_X97Y120_SLICE_X153Y120_A5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B5 = CLBLM_R_X97Y121_SLICE_X153Y121_DO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_B6 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C1 = CLBLM_R_X97Y120_SLICE_X153Y120_C5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C2 = CLBLM_L_X98Y121_SLICE_X155Y121_AQ;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C4 = CLBLL_L_X100Y121_SLICE_X157Y121_AQ;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C5 = CLBLM_R_X97Y120_SLICE_X153Y120_D5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_C6 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D1 = CLBLM_L_X94Y120_SLICE_X149Y120_B5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D3 = CLBLM_R_X95Y121_SLICE_X151Y121_DO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D4 = CLBLM_R_X97Y121_SLICE_X153Y121_A5Q;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D5 = CLBLM_R_X97Y123_SLICE_X153Y123_DO6;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y121_SLICE_X153Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A2 = CLBLM_R_X95Y121_SLICE_X150Y121_BO6;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A3 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A4 = CLBLM_R_X97Y122_SLICE_X152Y122_D5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A5 = CLBLM_R_X97Y122_SLICE_X153Y122_C5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_A6 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B2 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B3 = CLBLM_R_X97Y121_SLICE_X152Y121_AQ;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B4 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B5 = CLBLM_R_X97Y121_SLICE_X152Y121_C5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_B6 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C1 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C2 = CLBLM_R_X97Y121_SLICE_X152Y121_CQ;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C4 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C5 = CLBLM_R_X97Y122_SLICE_X152Y122_DQ;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_C6 = 1'b1;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D1 = CLBLM_R_X97Y121_SLICE_X152Y121_C5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D2 = CLBLM_R_X97Y121_SLICE_X152Y121_CQ;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D3 = CLBLM_R_X97Y122_SLICE_X152Y122_DQ;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D5 = CLBLM_R_X97Y121_SLICE_X152Y121_B5Q;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_D6 = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1 = 1'b0;
  assign CLBLM_R_X97Y121_SLICE_X152Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign LIOI3_X0Y227_OLOGIC_X0Y228_D1 = 1'b0;
  assign LIOI3_X0Y227_OLOGIC_X0Y228_T1 = 1'b1;
  assign LIOI3_X0Y227_OLOGIC_X0Y227_D1 = 1'b0;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = 1'b0;
  assign LIOI3_X0Y227_OLOGIC_X0Y227_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b0;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = 1'b0;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = 1'b0;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = 1'b0;
  assign LIOB33_X0Y171_IOB_X0Y172_O = 1'b0;
  assign LIOB33_X0Y171_IOB_X0Y171_O = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign LIOB33_X0Y171_IOB_X0Y172_T = 1'b1;
  assign LIOB33_X0Y171_IOB_X0Y171_T = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A2 = CLBLM_L_X98Y123_SLICE_X154Y123_CQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A3 = CLBLM_R_X97Y122_SLICE_X153Y122_AQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A4 = CLBLM_L_X98Y122_SLICE_X154Y122_B5Q;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A5 = CLBLM_R_X97Y122_SLICE_X152Y122_CQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_A6 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B2 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B3 = CLBLM_L_X98Y122_SLICE_X155Y122_B5Q;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B4 = CLBLL_L_X100Y123_SLICE_X156Y123_AQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B5 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_B6 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C1 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C2 = CLBLM_R_X97Y122_SLICE_X153Y122_CQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C4 = CLBLM_R_X97Y122_SLICE_X153Y122_BQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C5 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_C6 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D1 = CLBLM_R_X97Y122_SLICE_X153Y122_C5Q;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D2 = CLBLM_R_X97Y122_SLICE_X153Y122_CQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D3 = CLBLL_L_X100Y123_SLICE_X156Y123_AQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D4 = CLBLM_R_X97Y122_SLICE_X153Y122_BQ;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_D6 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X153Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A2 = CLBLM_R_X97Y122_SLICE_X152Y122_A5Q;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A3 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A4 = CLBLM_L_X98Y122_SLICE_X154Y122_AQ;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A5 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_A6 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B2 = CLBLM_R_X93Y122_SLICE_X146Y122_BO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B3 = CLBLM_L_X98Y121_SLICE_X154Y121_BO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B5 = CLBLM_R_X97Y122_SLICE_X152Y122_A5Q;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_B6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C1 = CLBLM_L_X98Y122_SLICE_X154Y122_AQ;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C5 = CLBLM_R_X93Y123_SLICE_X146Y123_CO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_C6 = CLBLM_R_X97Y122_SLICE_X153Y122_AO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D1 = CLBLM_R_X95Y121_SLICE_X150Y121_CO6;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D2 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D3 = CLBLM_R_X97Y122_SLICE_X153Y122_B5Q;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D4 = CLBLM_R_X95Y122_SLICE_X150Y122_A5Q;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_D6 = 1'b1;
  assign CLBLM_R_X97Y122_SLICE_X152Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1 = CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B5 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B6 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y174_O = 1'b0;
  assign LIOB33_X0Y173_IOB_X0Y173_O = 1'b0;
  assign LIOB33_X0Y173_IOB_X0Y174_T = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y173_T = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A2 = CLBLM_R_X95Y122_SLICE_X151Y122_AO6;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A3 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A4 = CLBLM_R_X97Y121_SLICE_X153Y121_B5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A5 = CLBLM_R_X97Y123_SLICE_X153Y123_B5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_A6 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B2 = CLBLM_R_X97Y123_SLICE_X153Y123_BQ;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B3 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B4 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B5 = CLBLM_L_X98Y124_SLICE_X154Y124_AQ;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_B6 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C1 = CLBLM_L_X98Y123_SLICE_X154Y123_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C2 = CLBLM_R_X97Y123_SLICE_X153Y123_CQ;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_AX = CLBLM_L_X92Y131_SLICE_X145Y131_BO5;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C4 = CLBLM_R_X97Y121_SLICE_X153Y121_C5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C5 = CLBLM_L_X98Y123_SLICE_X155Y123_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_C6 = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_D1 = 1'b0;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B1 = CLBLM_L_X92Y131_SLICE_X144Y131_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D1 = CLBLM_L_X98Y124_SLICE_X154Y124_AQ;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B2 = CLBLM_L_X92Y131_SLICE_X145Y131_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D3 = CLBLM_R_X97Y123_SLICE_X153Y123_BQ;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D4 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D5 = CLBLM_R_X97Y123_SLICE_X153Y123_B5Q;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_D6 = CLBLL_L_X100Y124_SLICE_X157Y124_BQ;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B3 = CLBLM_L_X92Y131_SLICE_X145Y131_AQ;
  assign CLBLM_R_X97Y123_SLICE_X153Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A2 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A3 = CLBLM_R_X97Y123_SLICE_X153Y123_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A4 = CLBLM_R_X97Y125_SLICE_X153Y125_A5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A5 = CLBLM_R_X95Y123_SLICE_X151Y123_CO6;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_A6 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B2 = CLBLM_R_X97Y123_SLICE_X152Y123_BQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B3 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B4 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B5 = CLBLM_R_X97Y124_SLICE_X152Y124_BQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_B6 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C1 = CLBLM_R_X97Y122_SLICE_X153Y122_AQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C2 = CLBLM_R_X97Y123_SLICE_X152Y123_CQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C4 = CLBLM_L_X98Y121_SLICE_X154Y121_BQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C5 = CLBLM_R_X97Y123_SLICE_X153Y123_C5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_C6 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D1 = CLBLM_L_X98Y125_SLICE_X154Y125_AQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D2 = CLBLM_R_X97Y124_SLICE_X152Y124_BQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D3 = 1'b1;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D4 = CLBLM_R_X97Y123_SLICE_X152Y123_BQ;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D5 = CLBLM_R_X97Y123_SLICE_X152Y123_B5Q;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y123_SLICE_X152Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1 = 1'b0;
  assign LIOB33_X0Y175_IOB_X0Y176_O = 1'b0;
  assign LIOB33_X0Y175_IOB_X0Y175_O = 1'b0;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_T = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y175_T = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1 = 1'b0;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D5 = 1'b1;
  assign LIOI3_X0Y229_OLOGIC_X0Y230_D1 = 1'b0;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y229_OLOGIC_X0Y230_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1 = 1'b1;
  assign LIOI3_X0Y229_OLOGIC_X0Y229_D1 = 1'b0;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = 1'b0;
  assign LIOI3_X0Y229_OLOGIC_X0Y229_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b0;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A1 = CLBLM_R_X97Y123_SLICE_X152Y123_DO6;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A2 = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A5 = CLBLM_R_X97Y124_SLICE_X152Y124_AQ;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_A6 = CLBLM_R_X95Y122_SLICE_X150Y122_A5Q;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = 1'b0;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B2 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B3 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B4 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B5 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_B6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = 1'b0;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b0;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C2 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C3 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C4 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C5 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D2 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D3 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D4 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D5 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X153Y124_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = 1'b0;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A2 = CLBLM_R_X97Y124_SLICE_X152Y124_A5Q;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A3 = CLBLM_R_X95Y125_SLICE_X150Y125_AQ;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A4 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A5 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B2 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B3 = CLBLM_L_X98Y125_SLICE_X154Y125_AQ;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B4 = CLBLM_R_X95Y124_SLICE_X151Y124_CQ;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B5 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_B6 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C1 = CLBLM_R_X97Y124_SLICE_X152Y124_A5Q;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C2 = CLBLM_L_X94Y124_SLICE_X149Y124_CO6;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C3 = CLBLM_R_X95Y124_SLICE_X150Y124_B5Q;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C4 = CLBLM_L_X98Y127_SLICE_X155Y127_CO6;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOB33_X105Y179_IOB_X1Y180_T = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D1 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D2 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D3 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D4 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D5 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_D6 = 1'b1;
  assign CLBLM_R_X97Y124_SLICE_X152Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y179_IOB_X1Y179_T = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A1 = CLBLM_R_X95Y113_SLICE_X150Y113_B5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A2 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A3 = CLBLM_R_X93Y114_SLICE_X147Y114_A5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A5 = CLBLM_L_X94Y111_SLICE_X149Y111_CO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_A6 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D2 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B1 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B3 = CLBLM_L_X94Y111_SLICE_X149Y111_AQ;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B4 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B5 = CLBLM_L_X94Y111_SLICE_X149Y111_BQ;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_B6 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D3 = CLBLM_L_X92Y112_SLICE_X145Y112_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D4 = CLBLM_R_X93Y112_SLICE_X146Y112_BQ;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C1 = CLBLM_L_X94Y112_SLICE_X149Y112_A5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C2 = CLBLM_R_X97Y111_SLICE_X152Y111_A5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C3 = CLBLM_R_X93Y112_SLICE_X147Y112_DO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C5 = CLBLM_L_X94Y111_SLICE_X149Y111_DO6;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D1 = CLBLM_L_X94Y111_SLICE_X149Y111_BQ;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D2 = CLBLM_R_X95Y111_SLICE_X150Y111_B5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D3 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D4 = CLBLM_L_X94Y111_SLICE_X149Y111_AQ;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D5 = CLBLM_L_X94Y111_SLICE_X149Y111_B5Q;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = 1'b0;
  assign LIOB33_X0Y177_IOB_X0Y177_O = 1'b0;
  assign CLBLM_L_X94Y111_SLICE_X149Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B1 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A1 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A2 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A3 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A4 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A5 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_A6 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B2 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y177_T = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_T = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B1 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B2 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B3 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B4 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B5 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_B6 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C1 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C2 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C3 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C4 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C5 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_C6 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D1 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D2 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D3 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D4 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D5 = 1'b1;
  assign CLBLM_L_X94Y111_SLICE_X148Y111_D6 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A2 = CLBLM_L_X98Y126_SLICE_X154Y126_BQ;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A3 = CLBLM_R_X97Y125_SLICE_X152Y125_B5Q;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A4 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C6 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A5 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_A6 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B2 = CLBLM_R_X97Y125_SLICE_X153Y125_BQ;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B3 = CLBLM_R_X97Y125_SLICE_X153Y125_AQ;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B4 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B5 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_B6 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C2 = CLBLM_R_X97Y125_SLICE_X152Y125_CO6;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C3 = CLBLL_L_X100Y126_SLICE_X156Y126_CO6;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C4 = CLBLM_R_X97Y123_SLICE_X152Y123_A5Q;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_C6 = CLBLM_L_X98Y125_SLICE_X154Y125_B5Q;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D2 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D3 = CLBLM_R_X97Y125_SLICE_X153Y125_BQ;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D4 = CLBLM_R_X97Y125_SLICE_X153Y125_AQ;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D5 = CLBLM_R_X97Y125_SLICE_X153Y125_B5Q;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_D6 = CLBLM_L_X98Y126_SLICE_X154Y126_BQ;
  assign CLBLM_R_X97Y125_SLICE_X153Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A2 = CLBLM_R_X95Y125_SLICE_X151Y125_BO6;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A3 = CLBLM_R_X97Y125_SLICE_X153Y125_B5Q;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A4 = CLBLM_R_X97Y123_SLICE_X152Y123_A5Q;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A5 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_A6 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B2 = CLBLM_R_X97Y125_SLICE_X152Y125_BQ;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B3 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B4 = CLBLM_L_X98Y125_SLICE_X154Y125_CQ;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B5 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_B6 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C2 = CLBLM_R_X97Y125_SLICE_X153Y125_A5Q;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C3 = CLBLM_R_X97Y125_SLICE_X152Y125_BQ;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C4 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C5 = CLBLM_R_X97Y125_SLICE_X152Y125_B5Q;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_C6 = CLBLM_L_X98Y125_SLICE_X154Y125_CQ;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D1 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D2 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D3 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D4 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D5 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_D6 = 1'b1;
  assign CLBLM_R_X97Y125_SLICE_X152Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A1 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A3 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A4 = CLBLM_R_X95Y113_SLICE_X151Y113_AQ;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A5 = CLBLM_L_X94Y112_SLICE_X149Y112_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_A6 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B2 = CLBLM_R_X93Y112_SLICE_X147Y112_C5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B3 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B4 = CLBLM_L_X94Y111_SLICE_X149Y111_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B5 = CLBLM_L_X94Y112_SLICE_X149Y112_CO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_B6 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = 1'b0;
  assign LIOB33_X0Y179_IOB_X0Y180_O = 1'b0;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C3 = CLBLM_L_X94Y114_SLICE_X148Y114_CO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C4 = CLBLM_R_X95Y111_SLICE_X150Y111_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C5 = CLBLM_R_X95Y111_SLICE_X150Y111_DO6;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_C6 = CLBLM_L_X94Y112_SLICE_X149Y112_AQ;
  assign LIOB33_X0Y179_IOB_X0Y179_T = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_T = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D1 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D2 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D3 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D4 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D5 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_D6 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X149Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A1 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A2 = CLBLM_L_X94Y112_SLICE_X148Y112_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A3 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A5 = CLBLM_L_X94Y112_SLICE_X149Y112_AQ;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y77_IOB_X1Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B1 = CLBLM_L_X94Y112_SLICE_X148Y112_DO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B2 = CLBLM_R_X93Y113_SLICE_X147Y113_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B3 = CLBLM_L_X94Y112_SLICE_X149Y112_B5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B5 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_B6 = 1'b1;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C1 = CLBLM_R_X93Y112_SLICE_X146Y112_DO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C2 = CLBLM_R_X95Y112_SLICE_X150Y112_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C3 = CLBLM_L_X94Y112_SLICE_X148Y112_AQ;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C4 = CLBLM_R_X93Y111_SLICE_X147Y111_CO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D1 = CLBLM_L_X94Y112_SLICE_X148Y112_A5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D2 = CLBLM_R_X95Y112_SLICE_X150Y112_B5Q;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D3 = CLBLM_R_X93Y113_SLICE_X147Y113_DO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D5 = CLBLM_R_X93Y112_SLICE_X146Y112_CO6;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y112_SLICE_X148Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b0;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A2 = CLBLM_R_X97Y126_SLICE_X153Y126_BQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A3 = CLBLM_R_X97Y126_SLICE_X153Y126_AQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A4 = CLBLM_R_X97Y127_SLICE_X153Y127_BQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A5 = CLBLM_R_X97Y126_SLICE_X153Y126_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_A6 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B2 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B3 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B4 = CLBLM_R_X97Y127_SLICE_X153Y127_BQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B5 = CLBLM_R_X97Y126_SLICE_X153Y126_BQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_B6 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C1 = CLBLM_R_X97Y128_SLICE_X152Y128_AQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C2 = CLBLM_R_X97Y126_SLICE_X153Y126_CQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C3 = CLBLM_L_X94Y127_SLICE_X149Y127_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C4 = CLBLM_L_X94Y125_SLICE_X149Y125_A5Q;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_C6 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D1 = CLBLM_R_X97Y126_SLICE_X153Y126_BQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D2 = CLBLM_R_X97Y126_SLICE_X153Y126_CQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D4 = CLBLM_R_X97Y126_SLICE_X153Y126_AQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D5 = CLBLM_R_X97Y126_SLICE_X153Y126_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_D6 = CLBLM_R_X97Y127_SLICE_X153Y127_BQ;
  assign CLBLM_R_X97Y126_SLICE_X153Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A2 = CLBLM_R_X97Y127_SLICE_X152Y127_A5Q;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A3 = CLBLM_R_X97Y125_SLICE_X152Y125_A5Q;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A4 = CLBLM_R_X95Y126_SLICE_X151Y126_BO6;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A5 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_A6 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B2 = CLBLM_R_X97Y126_SLICE_X152Y126_BQ;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B3 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B4 = CLBLM_L_X98Y127_SLICE_X154Y127_BQ;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B5 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_B6 = 1'b1;
  assign LIOI3_X0Y233_OLOGIC_X0Y234_D1 = 1'b0;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C2 = CLBLM_R_X97Y127_SLICE_X152Y127_A5Q;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C3 = CLBLM_R_X97Y126_SLICE_X152Y126_BQ;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C4 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C5 = CLBLM_R_X97Y126_SLICE_X152Y126_B5Q;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_C6 = CLBLM_L_X98Y127_SLICE_X154Y127_BQ;
  assign LIOI3_X0Y233_OLOGIC_X0Y234_T1 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D1 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D2 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D3 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D4 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D5 = 1'b1;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_D6 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_O = 1'b0;
  assign LIOB33_X0Y181_IOB_X0Y182_O = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = 1'b0;
  assign CLBLM_R_X97Y126_SLICE_X152Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y233_OLOGIC_X0Y233_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_T = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_T = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A2 = CLBLM_R_X95Y114_SLICE_X150Y114_BQ;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A3 = CLBLM_L_X94Y113_SLICE_X149Y113_AQ;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A5 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_A6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B1 = CLBLM_L_X94Y116_SLICE_X149Y116_BQ;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B3 = CLBLM_R_X95Y113_SLICE_X150Y113_B5Q;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B5 = CLBLM_L_X94Y115_SLICE_X149Y115_DO6;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_B6 = CLBLM_L_X94Y113_SLICE_X149Y113_CO6;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = 1'b0;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C2 = CLBLM_R_X95Y114_SLICE_X150Y114_BQ;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C4 = CLBLM_L_X94Y113_SLICE_X149Y113_A5Q;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C5 = CLBLM_L_X94Y113_SLICE_X149Y113_AQ;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_C6 = CLBLM_L_X94Y114_SLICE_X149Y114_BQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b0;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D2 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D3 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D4 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D5 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X149Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A1 = CLBLM_L_X94Y114_SLICE_X149Y114_CO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A2 = CLBLM_L_X92Y113_SLICE_X144Y113_A5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A3 = CLBLM_R_X95Y112_SLICE_X150Y112_A5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A5 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B1 = CLBLM_L_X94Y113_SLICE_X148Y113_B5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B3 = CLBLM_L_X94Y114_SLICE_X148Y114_AQ;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B4 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B5 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_B6 = 1'b1;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C2 = CLBLM_L_X94Y114_SLICE_X148Y114_CO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C4 = CLBLM_L_X94Y112_SLICE_X148Y112_B5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C5 = CLBLM_L_X94Y113_SLICE_X148Y113_B5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_C6 = CLBLM_L_X94Y116_SLICE_X148Y116_DO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D1 = CLBLM_L_X94Y114_SLICE_X148Y114_AQ;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D2 = CLBLM_R_X93Y112_SLICE_X147Y112_DO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D5 = CLBLM_L_X94Y112_SLICE_X149Y112_B5Q;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_D6 = CLBLM_L_X94Y117_SLICE_X148Y117_DO6;
  assign CLBLM_L_X94Y113_SLICE_X148Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A2 = CLBLM_R_X97Y126_SLICE_X152Y126_A5Q;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A3 = CLBLM_R_X97Y127_SLICE_X152Y127_CO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A4 = CLBLM_R_X97Y127_SLICE_X152Y127_B5Q;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A5 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_A6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = 1'b0;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLL_L_X102Y123_SLICE_X160Y123_CO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B1 = CLBLM_R_X101Y127_SLICE_X159Y127_BO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B3 = CLBLM_R_X97Y126_SLICE_X153Y126_AO6;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B5 = CLBLM_R_X97Y129_SLICE_X152Y129_AQ;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C1 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C2 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C3 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C4 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C5 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_C6 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D1 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D2 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D3 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D4 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D5 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_D6 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X153Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A2 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A3 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A4 = CLBLM_R_X97Y126_SLICE_X152Y126_B5Q;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A5 = CLBLM_L_X98Y127_SLICE_X155Y127_AQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_A6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y183_O = 1'b0;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B2 = CLBLM_R_X97Y127_SLICE_X152Y127_BQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B3 = CLBLM_R_X97Y127_SLICE_X152Y127_AQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B4 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B5 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_B6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y184_O = 1'b0;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_T1 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y184_T = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C1 = CLBLM_R_X95Y124_SLICE_X150Y124_C5Q;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C2 = CLBLM_R_X95Y125_SLICE_X151Y125_CO6;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C3 = CLBLM_R_X95Y126_SLICE_X151Y126_AQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C5 = CLBLM_L_X98Y128_SLICE_X154Y128_DO6;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y183_IOB_X0Y183_T = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D1 = CLBLM_L_X98Y127_SLICE_X155Y127_AQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D2 = CLBLM_R_X97Y127_SLICE_X152Y127_AQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D3 = CLBLM_R_X97Y127_SLICE_X152Y127_BQ;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D4 = 1'b1;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D5 = CLBLM_R_X97Y127_SLICE_X152Y127_B5Q;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y127_SLICE_X152Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A1 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A2 = CLBLM_L_X94Y114_SLICE_X149Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A4 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A5 = CLBLM_R_X95Y113_SLICE_X150Y113_AQ;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_A6 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B1 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B2 = CLBLM_L_X94Y113_SLICE_X149Y113_BO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B4 = CLBLM_L_X94Y115_SLICE_X149Y115_CO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B5 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_D1 = 1'b0;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C1 = CLBLM_L_X92Y113_SLICE_X144Y113_CO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C2 = CLBLM_R_X95Y116_SLICE_X150Y116_CO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C4 = CLBLM_L_X94Y114_SLICE_X149Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C5 = CLBLM_L_X98Y114_SLICE_X154Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D1 = CLBLM_L_X94Y111_SLICE_X149Y111_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D2 = CLBLM_L_X94Y114_SLICE_X148Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D3 = CLBLM_R_X93Y114_SLICE_X147Y114_CO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D4 = CLBLM_L_X94Y117_SLICE_X149Y117_DO6;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y114_SLICE_X149Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A1 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A2 = CLBLM_L_X94Y114_SLICE_X148Y114_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A3 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A4 = CLBLM_L_X94Y116_SLICE_X149Y116_BQ;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_A6 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B1 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B2 = CLBLM_L_X94Y114_SLICE_X148Y114_BQ;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B3 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B4 = CLBLM_L_X94Y115_SLICE_X148Y115_BQ;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_B6 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C1 = CLBLM_L_X94Y114_SLICE_X148Y114_BQ;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C2 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C4 = CLBLM_R_X93Y113_SLICE_X147Y113_A5Q;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C5 = CLBLM_L_X94Y114_SLICE_X148Y114_B5Q;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_C6 = CLBLM_L_X94Y115_SLICE_X148Y115_BQ;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y219_T1 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D1 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D2 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D3 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D4 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D5 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_D6 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B4 = 1'b1;
  assign CLBLM_L_X94Y114_SLICE_X148Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B3 = CLBLL_L_X102Y119_SLICE_X160Y119_AQ;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B4 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B5 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B6 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A1 = CLBLM_R_X97Y129_SLICE_X152Y129_A5Q;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A2 = CLBLL_L_X102Y128_SLICE_X161Y128_DO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A3 = CLBLM_R_X93Y132_SLICE_X146Y132_AQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A4 = CLBLM_R_X97Y128_SLICE_X153Y128_BO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A4 = CLBLM_L_X92Y132_SLICE_X145Y132_BO6;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_AX = CLBLM_R_X97Y128_SLICE_X153Y128_BO5;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B2 = CLBLM_R_X97Y128_SLICE_X153Y128_A5Q;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B3 = CLBLM_R_X97Y128_SLICE_X153Y128_AQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B4 = CLBLM_R_X97Y128_SLICE_X153Y128_CQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B5 = CLBLM_R_X97Y128_SLICE_X153Y128_C5Q;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_B6 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C1 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C2 = CLBLM_R_X97Y128_SLICE_X153Y128_CQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C3 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C5 = CLBLM_R_X97Y128_SLICE_X153Y128_AQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_C6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = 1'b0;
  assign LIOB33_X0Y185_IOB_X0Y185_O = 1'b0;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D1 = CLBLM_R_X97Y128_SLICE_X153Y128_C5Q;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D3 = CLBLM_R_X97Y128_SLICE_X152Y128_AQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D4 = CLBLM_R_X97Y128_SLICE_X153Y128_A5Q;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D5 = CLBLM_R_X97Y128_SLICE_X153Y128_AQ;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_D6 = CLBLM_R_X97Y128_SLICE_X153Y128_CQ;
  assign LIOB33_X0Y185_IOB_X0Y185_T = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_T = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X153Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D2 = CLBLL_L_X102Y119_SLICE_X160Y119_AQ;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A2 = CLBLM_L_X94Y128_SLICE_X149Y128_A5Q;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A3 = CLBLM_R_X97Y129_SLICE_X152Y129_CQ;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A4 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A5 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A4 = CLBLM_L_X98Y116_SLICE_X155Y116_CO6;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_A6 = CLBLM_R_X95Y124_SLICE_X150Y124_C5Q;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D4 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B1 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B2 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B3 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B4 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B5 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_B6 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C1 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C2 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C3 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C4 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C5 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_C6 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D1 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D2 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D3 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D4 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D5 = 1'b1;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_D6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B2 = CLBLL_L_X100Y117_SLICE_X156Y117_BQ;
  assign CLBLM_R_X97Y128_SLICE_X152Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A2 = CLBLM_R_X95Y121_SLICE_X150Y121_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A3 = CLBLM_L_X94Y116_SLICE_X149Y116_C5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A4 = CLBLM_L_X94Y114_SLICE_X149Y114_DO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A5 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_A6 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B2 = CLBLM_L_X94Y115_SLICE_X149Y115_BQ;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B3 = CLBLM_L_X94Y114_SLICE_X149Y114_B5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B4 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B5 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_B6 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C2 = CLBLM_L_X94Y117_SLICE_X149Y117_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C4 = CLBLM_L_X94Y115_SLICE_X149Y115_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C5 = CLBLM_L_X94Y115_SLICE_X149Y115_DO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_C6 = CLBLM_R_X101Y121_SLICE_X159Y121_DO6;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C1 = CLBLL_L_X100Y117_SLICE_X157Y117_AQ;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D1 = CLBLM_L_X94Y116_SLICE_X149Y116_C5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D2 = CLBLM_L_X94Y114_SLICE_X149Y114_B5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D3 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D4 = CLBLM_L_X94Y115_SLICE_X149Y115_BQ;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D5 = CLBLM_L_X94Y115_SLICE_X149Y115_B5Q;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y115_SLICE_X149Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C4 = CLBLL_L_X102Y116_SLICE_X160Y116_C5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A2 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A3 = CLBLM_L_X94Y115_SLICE_X148Y115_AQ;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A4 = CLBLM_R_X95Y115_SLICE_X150Y115_AQ;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A5 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_A6 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B2 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B3 = CLBLM_L_X94Y117_SLICE_X148Y117_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B4 = CLBLM_L_X94Y113_SLICE_X148Y113_CO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B5 = CLBLM_L_X94Y115_SLICE_X148Y115_C5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_B6 = 1'b1;
  assign LIOI3_X0Y235_OLOGIC_X0Y236_D1 = 1'b0;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C1 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C2 = CLBLM_L_X94Y115_SLICE_X149Y115_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C3 = CLBLM_L_X94Y113_SLICE_X148Y113_DO6;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C5 = CLBLM_L_X94Y117_SLICE_X149Y117_B5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_C6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y235_OLOGIC_X0Y236_T1 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D1 = CLBLM_R_X95Y115_SLICE_X150Y115_AQ;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D2 = 1'b1;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D3 = CLBLM_L_X94Y115_SLICE_X148Y115_AQ;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D4 = CLBLM_L_X94Y115_SLICE_X148Y115_A5Q;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_D6 = CLBLM_R_X93Y115_SLICE_X147Y115_AQ;
  assign LIOI3_X0Y235_OLOGIC_X0Y235_D1 = 1'b0;
  assign CLBLM_L_X94Y115_SLICE_X148Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = 1'b0;
  assign LIOI3_X0Y235_OLOGIC_X0Y235_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = 1'b0;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b0;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D3 = CLBLM_R_X101Y126_SLICE_X159Y126_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = 1'b0;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D4 = CLBLM_R_X103Y126_SLICE_X162Y126_BQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D5 = CLBLM_R_X103Y126_SLICE_X162Y126_B5Q;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B6 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y187_IOB_X0Y188_O = 1'b0;
  assign LIOB33_X0Y187_IOB_X0Y187_O = 1'b0;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A1 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A2 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A3 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A4 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_A6 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_T = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y187_T = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B1 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B2 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B3 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B4 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_B6 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C1 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C2 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C3 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C4 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_C6 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D1 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D2 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D3 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D4 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X153Y129_D6 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A1 = CLBLM_L_X98Y133_SLICE_X154Y133_AQ;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A2 = CLBLM_R_X97Y129_SLICE_X152Y129_A5Q;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A3 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_A6 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B1 = CLBLM_R_X97Y131_SLICE_X153Y131_CQ;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B2 = CLBLM_L_X94Y129_SLICE_X148Y129_AQ;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B3 = CLBLM_R_X95Y124_SLICE_X150Y124_C5Q;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B5 = CLBLM_R_X95Y129_SLICE_X150Y129_A5Q;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_B6 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C1 = CLBLM_R_X97Y132_SLICE_X153Y132_C5Q;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C2 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C3 = CLBLM_R_X95Y128_SLICE_X150Y128_AQ;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C4 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_C6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D1 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D2 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D3 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D4 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D5 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_D6 = 1'b1;
  assign CLBLM_R_X97Y129_SLICE_X152Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A2 = CLBLM_R_X97Y115_SLICE_X152Y115_A5Q;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A3 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A4 = CLBLM_R_X93Y116_SLICE_X146Y116_A5Q;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A5 = CLBLM_L_X98Y117_SLICE_X155Y117_CO6;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_A6 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B2 = CLBLM_L_X94Y120_SLICE_X148Y120_AQ;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B3 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B4 = CLBLM_L_X94Y116_SLICE_X149Y116_B5Q;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B5 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_B6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D4 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C1 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C2 = CLBLM_L_X94Y115_SLICE_X149Y115_B5Q;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C4 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C5 = CLBLM_R_X95Y117_SLICE_X150Y117_AQ;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_C6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D5 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D1 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D2 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D3 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D4 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D5 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_D6 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X149Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A2 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A3 = CLBLM_L_X94Y116_SLICE_X148Y116_AQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A4 = CLBLM_L_X94Y120_SLICE_X149Y120_BQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A5 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_A6 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B2 = CLBLM_L_X94Y116_SLICE_X148Y116_BQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B3 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B4 = CLBLM_L_X94Y117_SLICE_X148Y117_AQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B5 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_B6 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C1 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C2 = CLBLM_L_X94Y116_SLICE_X148Y116_AQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C4 = CLBLM_L_X94Y116_SLICE_X148Y116_A5Q;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C5 = CLBLM_R_X93Y116_SLICE_X147Y116_A5Q;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_C6 = CLBLM_L_X94Y120_SLICE_X149Y120_BQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D1 = CLBLM_R_X95Y118_SLICE_X150Y118_AQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D2 = 1'b1;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D4 = CLBLM_L_X94Y116_SLICE_X148Y116_BQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D5 = CLBLM_L_X94Y116_SLICE_X148Y116_B5Q;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_D6 = CLBLM_L_X94Y117_SLICE_X148Y117_AQ;
  assign CLBLM_L_X94Y116_SLICE_X148Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y189_IOB_X0Y190_O = 1'b0;
  assign LIOB33_X0Y189_IOB_X0Y189_O = 1'b0;
  assign LIOB33_X0Y189_IOB_X0Y190_T = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y189_T = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A2 = CLBLM_R_X95Y129_SLICE_X151Y129_B5Q;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A3 = CLBLM_R_X97Y130_SLICE_X153Y130_AQ;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A4 = CLBLM_R_X97Y129_SLICE_X152Y129_BQ;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A5 = CLBLM_R_X95Y130_SLICE_X151Y130_A5Q;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_A6 = 1'b1;
  assign LIOB33_X0Y87_IOB_X0Y88_O = 1'b0;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B1 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B2 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B3 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B4 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B5 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_B6 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C1 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C2 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C3 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C4 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C5 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_C6 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D1 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D2 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D3 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D4 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D5 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_D6 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X153Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A1 = CLBLM_R_X97Y130_SLICE_X152Y130_B5Q;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A2 = CLBLM_R_X97Y130_SLICE_X152Y130_BQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A3 = CLBLM_R_X97Y130_SLICE_X152Y130_AQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A4 = CLBLM_L_X98Y131_SLICE_X155Y131_BQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_A6 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B2 = CLBLM_R_X97Y130_SLICE_X152Y130_BQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B3 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B4 = CLBLM_L_X98Y131_SLICE_X155Y131_BQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B5 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_B6 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C1 = CLBLM_R_X97Y130_SLICE_X152Y130_BQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C2 = CLBLM_R_X97Y130_SLICE_X152Y130_AQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C3 = CLBLM_R_X97Y129_SLICE_X152Y129_B5Q;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C5 = CLBLM_R_X97Y130_SLICE_X152Y130_B5Q;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_C6 = CLBLM_L_X98Y131_SLICE_X155Y131_BQ;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D1 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D2 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D3 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D4 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D5 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_D6 = 1'b1;
  assign CLBLM_R_X97Y130_SLICE_X152Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y135_IOB_X0Y136_O = 1'b0;
  assign LIOB33_X0Y135_IOB_X0Y135_O = 1'b0;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_T1 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A2 = CLBLM_L_X94Y117_SLICE_X149Y117_A5Q;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A3 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A4 = CLBLM_R_X95Y120_SLICE_X150Y120_AQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A5 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_A6 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B2 = CLBLM_L_X94Y117_SLICE_X149Y117_BQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B3 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B4 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B5 = CLBLM_L_X94Y116_SLICE_X149Y116_CQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_B6 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C1 = CLBLM_L_X94Y115_SLICE_X148Y115_C5Q;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C2 = CLBLM_L_X94Y117_SLICE_X149Y117_AQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C4 = CLBLM_R_X95Y117_SLICE_X150Y117_DO6;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C5 = CLBLM_L_X94Y117_SLICE_X149Y117_DO6;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D1 = CLBLM_L_X94Y117_SLICE_X149Y117_BQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D2 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D4 = CLBLM_R_X95Y117_SLICE_X150Y117_AQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D5 = CLBLM_L_X94Y117_SLICE_X149Y117_B5Q;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_D6 = CLBLM_L_X94Y116_SLICE_X149Y116_CQ;
  assign CLBLM_L_X94Y117_SLICE_X149Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A2 = CLBLM_R_X95Y118_SLICE_X150Y118_AQ;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A3 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A4 = CLBLM_L_X94Y117_SLICE_X148Y117_B5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A5 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_A6 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B2 = CLBLM_L_X94Y117_SLICE_X148Y117_BQ;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B3 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B4 = CLBLM_R_X95Y118_SLICE_X150Y118_BQ;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B5 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_B6 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C2 = CLBLM_L_X94Y118_SLICE_X148Y118_A5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C3 = CLBLM_L_X94Y115_SLICE_X148Y115_B5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C4 = CLBLM_R_X95Y118_SLICE_X151Y118_CO6;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C5 = CLBLM_L_X94Y117_SLICE_X148Y117_DO6;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D1 = CLBLM_L_X94Y117_SLICE_X148Y117_BQ;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D2 = 1'b1;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D4 = CLBLM_L_X94Y117_SLICE_X148Y117_A5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D5 = CLBLM_L_X94Y117_SLICE_X148Y117_B5Q;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_D6 = CLBLM_R_X95Y118_SLICE_X150Y118_BQ;
  assign CLBLM_L_X94Y117_SLICE_X148Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = 1'b0;
  assign RIOB33_X105Y165_IOB_X1Y165_O = 1'b0;
  assign LIOB33_X0Y191_IOB_X0Y192_O = 1'b0;
  assign LIOB33_X0Y191_IOB_X0Y191_O = 1'b0;
  assign LIOB33_X0Y191_IOB_X0Y192_T = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_T = 1'b1;
  assign LIOI3_X0Y239_OLOGIC_X0Y240_D1 = 1'b0;
  assign LIOI3_X0Y239_OLOGIC_X0Y240_T1 = 1'b1;
  assign LIOI3_X0Y239_OLOGIC_X0Y239_D1 = 1'b0;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A1 = CLBLM_R_X97Y132_SLICE_X153Y132_DO6;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A3 = CLBLM_R_X97Y131_SLICE_X152Y131_AO6;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A5 = CLBLM_R_X95Y131_SLICE_X150Y131_AQ;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = 1'b0;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B2 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B3 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B4 = CLBLM_L_X98Y132_SLICE_X155Y132_BQ;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B5 = CLBLM_R_X97Y131_SLICE_X153Y131_BQ;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_B6 = 1'b1;
  assign LIOI3_X0Y239_OLOGIC_X0Y239_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C1 = CLBLM_R_X97Y130_SLICE_X153Y130_A5Q;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C3 = CLBLM_R_X97Y129_SLICE_X152Y129_B5Q;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C4 = CLBLM_R_X95Y131_SLICE_X151Y131_A5Q;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C5 = CLBLM_R_X97Y131_SLICE_X152Y131_AQ;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_C6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = 1'b0;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = 1'b0;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D1 = CLBLM_R_X97Y131_SLICE_X153Y131_BQ;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D2 = CLBLM_R_X97Y131_SLICE_X153Y131_CQ;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D4 = CLBLM_L_X98Y131_SLICE_X155Y131_B5Q;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D5 = CLBLM_R_X97Y131_SLICE_X153Y131_B5Q;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A1 = CLBLM_R_X93Y112_SLICE_X147Y112_BQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A3 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A5 = CLBLM_R_X93Y112_SLICE_X146Y112_A5Q;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_A6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_D6 = CLBLM_L_X98Y132_SLICE_X155Y132_BQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B1 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B3 = CLBLM_R_X93Y111_SLICE_X147Y111_AQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B5 = CLBLM_R_X93Y111_SLICE_X147Y111_BQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_B6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A2 = CLBLM_R_X95Y131_SLICE_X151Y131_CQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A3 = CLBLM_R_X97Y131_SLICE_X152Y131_AQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A4 = CLBLM_R_X97Y131_SLICE_X152Y131_B5Q;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C2 = CLBLM_R_X93Y111_SLICE_X147Y111_AQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C3 = CLBLM_R_X93Y111_SLICE_X147Y111_BQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C4 = CLBLM_R_X93Y112_SLICE_X147Y112_BQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C5 = CLBLM_R_X93Y111_SLICE_X147Y111_B5Q;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_C6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B2 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B3 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B4 = CLBLM_R_X97Y132_SLICE_X152Y132_BQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B5 = CLBLM_R_X95Y131_SLICE_X151Y131_CQ;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D1 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D2 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D3 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D5 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_D6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C3 = CLBLM_R_X93Y131_SLICE_X147Y131_AQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C4 = CLBLM_R_X97Y132_SLICE_X152Y132_B5Q;
  assign CLBLM_R_X93Y111_SLICE_X147Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D1 = CLBLM_R_X97Y131_SLICE_X153Y131_AQ;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A1 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A2 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A3 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A5 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_A6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D3 = CLBLM_R_X97Y131_SLICE_X152Y131_AQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D4 = CLBLM_R_X95Y131_SLICE_X151Y131_CQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D5 = CLBLM_R_X97Y131_SLICE_X152Y131_B5Q;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B1 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B2 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B3 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B5 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_B6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C1 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C2 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C3 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C5 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_C6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A2 = CLBLM_L_X94Y119_SLICE_X148Y119_AQ;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A3 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A4 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A5 = CLBLM_L_X94Y118_SLICE_X149Y118_A5Q;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_A6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B1 = CLBLM_R_X95Y120_SLICE_X151Y120_CO6;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D1 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D2 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D3 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D4 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D5 = 1'b1;
  assign CLBLM_R_X93Y111_SLICE_X146Y111_D6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B5 = CLBLM_L_X94Y116_SLICE_X148Y116_CO6;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B6 = CLBLM_L_X94Y118_SLICE_X149Y118_A5Q;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C1 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C2 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C3 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C4 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C5 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_C6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D1 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D2 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D3 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D4 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D5 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_D6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A2 = CLBLM_L_X94Y118_SLICE_X148Y118_A5Q;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A3 = CLBLM_L_X94Y117_SLICE_X149Y117_AQ;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A4 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A5 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_A6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B1 = CLBLM_R_X97Y119_SLICE_X153Y119_DO6;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B2 = CLBLM_L_X94Y116_SLICE_X148Y116_DO6;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B3 = CLBLM_L_X94Y118_SLICE_X148Y118_AQ;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_B6 = CLBLM_R_X93Y115_SLICE_X147Y115_B5Q;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C1 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C2 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C3 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C4 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C5 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_C6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D1 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D2 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D3 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D4 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D5 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_D6 = 1'b1;
  assign CLBLM_L_X94Y118_SLICE_X148Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_SING_X0Y99_IOB_X0Y99_O = 1'b0;
  assign LIOB33_X0Y193_IOB_X0Y194_O = 1'b0;
  assign LIOB33_X0Y193_IOB_X0Y193_O = 1'b0;
  assign LIOB33_X0Y193_IOB_X0Y194_T = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_T = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A2 = CLBLM_L_X98Y133_SLICE_X155Y133_BQ;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A3 = CLBLM_R_X97Y132_SLICE_X153Y132_AQ;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A4 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A5 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_A6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B2 = CLBLM_R_X97Y132_SLICE_X153Y132_BQ;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B3 = CLBLM_R_X95Y132_SLICE_X151Y132_B5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B4 = CLBLM_R_X97Y132_SLICE_X152Y132_B5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B5 = CLBLM_R_X97Y131_SLICE_X153Y131_C5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_B6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C1 = CLBLM_R_X95Y132_SLICE_X150Y132_AQ;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C2 = CLBLM_R_X97Y132_SLICE_X153Y132_CQ;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C4 = CLBLM_R_X95Y130_SLICE_X150Y130_A5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C5 = CLBLM_R_X97Y132_SLICE_X153Y132_B5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_C6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D1 = CLBLM_L_X98Y132_SLICE_X155Y132_AQ;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D3 = CLBLM_R_X97Y131_SLICE_X153Y131_C5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D4 = CLBLM_R_X97Y132_SLICE_X153Y132_A5Q;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D5 = CLBLM_R_X97Y132_SLICE_X153Y132_AQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A1 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A2 = CLBLM_L_X94Y112_SLICE_X148Y112_AQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A3 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A5 = CLBLM_R_X93Y112_SLICE_X147Y112_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_A6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B1 = CLBLM_L_X94Y112_SLICE_X148Y112_B5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B2 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B3 = CLBLM_R_X93Y113_SLICE_X147Y113_B5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B4 = CLBLM_L_X94Y112_SLICE_X148Y112_CO6;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_B6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A2 = CLBLM_R_X97Y132_SLICE_X152Y132_A5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A3 = CLBLM_R_X95Y131_SLICE_X150Y131_AQ;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A4 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C2 = CLBLM_R_X93Y112_SLICE_X147Y112_CQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C3 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C4 = CLBLM_R_X93Y114_SLICE_X147Y114_AQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C5 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_C6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B2 = CLBLM_R_X97Y133_SLICE_X153Y133_DO6;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B5 = CLBLM_R_X97Y132_SLICE_X152Y132_A5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_BX = CLBLM_R_X97Y132_SLICE_X152Y132_CO5;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D1 = CLBLM_R_X93Y112_SLICE_X147Y112_C5Q;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D2 = CLBLM_R_X93Y112_SLICE_X147Y112_CQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D3 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D4 = CLBLM_R_X93Y114_SLICE_X147Y114_AQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_D6 = CLBLM_L_X94Y115_SLICE_X148Y115_CQ;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C4 = CLBLM_R_X97Y131_SLICE_X152Y131_BQ;
  assign CLBLM_R_X93Y112_SLICE_X147Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D1 = CLBLM_R_X97Y131_SLICE_X152Y131_BQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A1 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A3 = CLBLM_R_X93Y112_SLICE_X146Y112_AQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A4 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A5 = CLBLM_L_X94Y112_SLICE_X148Y112_BQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_A6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D3 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D4 = CLBLM_R_X95Y132_SLICE_X151Y132_CQ;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D5 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B1 = CLBLM_R_X93Y112_SLICE_X146Y112_BQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B3 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B4 = CLBLM_R_X93Y115_SLICE_X146Y115_BQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B5 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_B6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A1 = CLBLM_R_X95Y119_SLICE_X150Y119_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C2 = CLBLM_R_X93Y111_SLICE_X147Y111_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C3 = CLBLM_R_X93Y112_SLICE_X146Y112_AQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C4 = CLBLM_R_X93Y112_SLICE_X146Y112_A5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C5 = 1'b1;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_C6 = CLBLM_L_X94Y112_SLICE_X148Y112_BQ;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A3 = CLBLM_R_X95Y119_SLICE_X150Y119_C5Q;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A4 = CLBLM_L_X94Y119_SLICE_X148Y119_CO6;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A5 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_A6 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B1 = CLBLM_L_X94Y119_SLICE_X149Y119_BQ;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B3 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B4 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B5 = CLBLM_R_X95Y119_SLICE_X150Y119_AQ;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_B6 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C1 = CLBLM_R_X95Y119_SLICE_X150Y119_DO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C2 = CLBLM_L_X94Y119_SLICE_X148Y119_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C5 = CLBLM_L_X94Y119_SLICE_X149Y119_DO6;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_C6 = CLBLM_R_X93Y115_SLICE_X146Y115_B5Q;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D5 = CLBLM_R_X93Y112_SLICE_X146Y112_B5Q;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_D6 = CLBLM_R_X93Y115_SLICE_X146Y115_BQ;
  assign CLBLM_R_X93Y112_SLICE_X146Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D1 = CLBLM_R_X95Y119_SLICE_X150Y119_AQ;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D2 = CLBLM_R_X93Y118_SLICE_X147Y118_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D3 = CLBLM_L_X94Y119_SLICE_X149Y119_BQ;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D5 = CLBLM_L_X94Y119_SLICE_X149Y119_B5Q;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_D6 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X149Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A2 = CLBLM_L_X94Y119_SLICE_X148Y119_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A3 = CLBLM_L_X94Y118_SLICE_X148Y118_AQ;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A4 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A5 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_A6 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B1 = CLBLM_R_X93Y120_SLICE_X147Y120_DO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B4 = CLBLM_R_X97Y121_SLICE_X152Y121_DO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B5 = CLBLM_R_X93Y120_SLICE_X147Y120_C5Q;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_B6 = CLBLM_L_X94Y120_SLICE_X148Y120_AQ;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C1 = CLBLM_R_X95Y121_SLICE_X151Y121_DO6;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C2 = CLBLM_L_X94Y119_SLICE_X148Y119_AQ;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C3 = CLBLM_R_X93Y115_SLICE_X146Y115_A5Q;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_C6 = CLBLM_R_X93Y118_SLICE_X147Y118_CO6;
  assign LIOB33_X0Y195_IOB_X0Y196_O = 1'b0;
  assign LIOB33_X0Y195_IOB_X0Y195_O = 1'b0;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D1 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D2 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D3 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D4 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D5 = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_D6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y195_T = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_T = 1'b1;
  assign CLBLM_L_X94Y119_SLICE_X148Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A2 = CLBLM_L_X98Y133_SLICE_X155Y133_AQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A4 = CLBLM_R_X97Y133_SLICE_X153Y133_BO6;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A5 = CLBLM_R_X101Y136_SLICE_X159Y136_DO6;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_AX = CLBLM_R_X97Y133_SLICE_X153Y133_BO5;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B2 = CLBLM_R_X97Y133_SLICE_X153Y133_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B3 = CLBLM_R_X97Y133_SLICE_X153Y133_AQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B4 = CLBLM_R_X97Y133_SLICE_X153Y133_CQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B5 = CLBLM_R_X97Y133_SLICE_X153Y133_C5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_B6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C1 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C2 = CLBLM_R_X97Y133_SLICE_X153Y133_CQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C3 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C5 = CLBLM_R_X97Y133_SLICE_X153Y133_AQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_C6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D1 = CLBLM_R_X97Y133_SLICE_X153Y133_C5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D2 = CLBLM_R_X97Y133_SLICE_X153Y133_CQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D3 = CLBLM_R_X97Y132_SLICE_X153Y132_BQ;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D4 = CLBLM_R_X97Y133_SLICE_X153Y133_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D5 = CLBLM_R_X97Y133_SLICE_X153Y133_AQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A1 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A2 = CLBLM_R_X93Y115_SLICE_X147Y115_BQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A4 = CLBLM_L_X94Y114_SLICE_X148Y114_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A5 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_A6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A1 = CLBLM_L_X98Y133_SLICE_X154Y133_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B1 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B2 = CLBLM_R_X93Y113_SLICE_X147Y113_BQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B4 = CLBLM_R_X93Y113_SLICE_X147Y113_AQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B5 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_B6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A2 = CLBLM_R_X101Y135_SLICE_X158Y135_BO6;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A4 = CLBLM_R_X97Y133_SLICE_X152Y133_BO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C1 = CLBLM_L_X94Y113_SLICE_X148Y113_BQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C2 = CLBLM_R_X93Y112_SLICE_X147Y112_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C4 = CLBLM_L_X94Y119_SLICE_X149Y119_DO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C5 = CLBLM_R_X93Y113_SLICE_X147Y113_DO6;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_AX = CLBLM_R_X97Y133_SLICE_X152Y133_BO5;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B1 = CLBLM_R_X97Y133_SLICE_X152Y133_CQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B2 = CLBLM_R_X97Y133_SLICE_X152Y133_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B3 = CLBLM_R_X97Y133_SLICE_X152Y133_AQ;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B5 = CLBLM_R_X97Y133_SLICE_X152Y133_C5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D2 = CLBLM_R_X93Y113_SLICE_X147Y113_AQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D3 = CLBLM_R_X93Y113_SLICE_X147Y113_BQ;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D4 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D5 = CLBLM_R_X93Y113_SLICE_X147Y113_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_D6 = CLBLM_R_X93Y115_SLICE_X147Y115_BQ;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C3 = CLBLM_R_X97Y133_SLICE_X152Y133_AQ;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y113_SLICE_X147Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D1 = CLBLM_R_X97Y133_SLICE_X152Y133_C5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A1 = CLBLM_L_X92Y112_SLICE_X145Y112_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A2 = CLBLM_R_X93Y113_SLICE_X146Y113_CO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A3 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A4 = CLBLM_R_X93Y112_SLICE_X147Y112_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_A6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D2 = CLBLM_R_X97Y133_SLICE_X152Y133_CQ;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D4 = CLBLM_R_X97Y133_SLICE_X152Y133_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D5 = CLBLM_R_X97Y132_SLICE_X153Y132_C5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B1 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B2 = CLBLM_R_X93Y113_SLICE_X146Y113_BQ;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B3 = CLBLM_R_X93Y113_SLICE_X146Y113_AQ;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B5 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_B6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B6 = 1'b1;
  assign LIOI3_X0Y241_OLOGIC_X0Y242_T1 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A1 = CLBLM_L_X94Y120_SLICE_X149Y120_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C1 = CLBLM_L_X92Y112_SLICE_X145Y112_CO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C3 = CLBLM_L_X94Y113_SLICE_X148Y113_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C4 = CLBLM_R_X93Y112_SLICE_X147Y112_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C5 = CLBLM_R_X93Y113_SLICE_X146Y113_DO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A2 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A3 = CLBLM_R_X95Y120_SLICE_X151Y120_B5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A5 = CLBLM_L_X94Y120_SLICE_X149Y120_CO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_A6 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B1 = CLBLM_R_X95Y120_SLICE_X151Y120_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B2 = CLBLM_L_X94Y118_SLICE_X149Y118_BO6;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D2 = CLBLM_R_X93Y113_SLICE_X146Y113_AQ;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D3 = CLBLM_L_X92Y113_SLICE_X144Y113_A5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D4 = CLBLM_R_X93Y113_SLICE_X146Y113_BQ;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D5 = CLBLM_R_X93Y113_SLICE_X146Y113_B5Q;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_D6 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B5 = CLBLM_L_X94Y119_SLICE_X149Y119_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B6 = 1'b1;
  assign CLBLM_R_X93Y113_SLICE_X146Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C2 = CLBLM_R_X93Y116_SLICE_X147Y116_CO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C3 = CLBLM_L_X94Y118_SLICE_X149Y118_AQ;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C4 = CLBLM_R_X95Y123_SLICE_X150Y123_CO6;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_C6 = CLBLM_R_X93Y114_SLICE_X146Y114_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D1 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D2 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D3 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D4 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D5 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_D6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C6 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = 1'b0;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b0;
  assign LIOB33_X0Y197_IOB_X0Y197_O = 1'b0;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A1 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A2 = CLBLM_L_X94Y120_SLICE_X148Y120_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A3 = CLBLM_L_X92Y120_SLICE_X144Y120_AQ;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A5 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_A6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_T = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B1 = CLBLM_R_X95Y120_SLICE_X150Y120_B5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B3 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B4 = CLBLM_L_X94Y119_SLICE_X148Y119_BO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B5 = CLBLM_L_X94Y120_SLICE_X148Y120_C5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_B6 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_T = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_D1 = 1'b0;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C1 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C2 = CLBLM_R_X95Y122_SLICE_X150Y122_B5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C3 = CLBLM_R_X93Y124_SLICE_X147Y124_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C5 = CLBLM_L_X94Y120_SLICE_X148Y120_DO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_C6 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y237_T1 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D2 = CLBLM_R_X93Y120_SLICE_X147Y120_CQ;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D3 = CLBLM_R_X93Y120_SLICE_X146Y120_DO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D4 = CLBLM_L_X94Y120_SLICE_X148Y120_A5Q;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_D6 = CLBLM_R_X95Y120_SLICE_X150Y120_CO6;
  assign CLBLM_L_X94Y120_SLICE_X148Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C4 = CLBLM_L_X98Y112_SLICE_X154Y112_B5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C5 = CLBLM_R_X97Y112_SLICE_X152Y112_DO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C6 = CLBLM_R_X93Y111_SLICE_X147Y111_CO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D1 = CLBLM_R_X97Y111_SLICE_X153Y111_AQ;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D2 = CLBLM_L_X98Y111_SLICE_X155Y111_DO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D6 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D6 = CLBLM_L_X98Y112_SLICE_X155Y112_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A1 = CLBLM_R_X93Y114_SLICE_X147Y114_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A2 = CLBLM_L_X94Y115_SLICE_X148Y115_CQ;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A3 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A5 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_A6 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B1 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B2 = CLBLM_R_X93Y114_SLICE_X147Y114_BQ;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B3 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B5 = CLBLM_L_X94Y115_SLICE_X149Y115_AQ;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_B6 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C2 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C3 = CLBLM_R_X93Y114_SLICE_X147Y114_BQ;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C4 = CLBLM_R_X93Y114_SLICE_X147Y114_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C5 = CLBLM_R_X93Y114_SLICE_X147Y114_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_C6 = CLBLM_L_X94Y115_SLICE_X149Y115_AQ;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D1 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D2 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D3 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D4 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D5 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_D6 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X147Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y131_SLICE_X153Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A1 = CLBLM_R_X93Y116_SLICE_X147Y116_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A2 = CLBLM_L_X92Y114_SLICE_X144Y114_CO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A4 = CLBLM_R_X93Y114_SLICE_X146Y114_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A5 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_A6 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B1 = CLBLM_R_X93Y115_SLICE_X146Y115_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B2 = CLBLM_R_X93Y116_SLICE_X147Y116_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B4 = CLBLM_R_X93Y114_SLICE_X146Y114_DO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B5 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_B6 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A1 = CLBLM_L_X94Y118_SLICE_X149Y118_AQ;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C1 = CLBLM_L_X90Y113_SLICE_X143Y113_DO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C2 = CLBLM_R_X93Y112_SLICE_X147Y112_AQ;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C4 = CLBLM_L_X92Y113_SLICE_X144Y113_CO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C5 = CLBLM_R_X93Y115_SLICE_X147Y115_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A2 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A4 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A5 = CLBLM_L_X94Y121_SLICE_X149Y121_A5Q;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_A6 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B3 = CLBLM_L_X94Y121_SLICE_X149Y121_AQ;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B4 = CLBLM_R_X93Y119_SLICE_X146Y119_A5Q;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B5 = CLBLM_R_X93Y119_SLICE_X146Y119_DO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_B6 = CLBLM_R_X95Y126_SLICE_X150Y126_CO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C1 = CLBLM_L_X94Y121_SLICE_X149Y121_A5Q;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C2 = CLBLM_R_X93Y119_SLICE_X146Y119_B5Q;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C3 = CLBLM_R_X95Y123_SLICE_X151Y123_DO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_C6 = CLBLM_R_X93Y119_SLICE_X147Y119_CO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D1 = CLBLM_L_X90Y113_SLICE_X143Y113_DO6;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D2 = CLBLM_R_X93Y116_SLICE_X147Y116_CO6;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D5 = CLBLM_L_X92Y114_SLICE_X145Y114_A5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D6 = CLBLM_L_X90Y113_SLICE_X143Y113_A5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B6 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D1 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D2 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D3 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D4 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D5 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_D6 = 1'b1;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D5 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X149Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D6 = CLBLM_R_X101Y130_SLICE_X158Y130_C5Q;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A1 = CLBLM_L_X90Y121_SLICE_X143Y121_DO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A4 = CLBLM_L_X94Y121_SLICE_X148Y121_BO6;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_A6 = CLBLM_L_X92Y119_SLICE_X145Y119_AQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_AX = CLBLM_L_X94Y121_SLICE_X148Y121_BO5;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B1 = CLBLM_L_X94Y121_SLICE_X148Y121_CQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B2 = CLBLM_L_X94Y121_SLICE_X148Y121_A5Q;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B3 = CLBLM_L_X94Y121_SLICE_X148Y121_AQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B4 = CLBLM_R_X93Y121_SLICE_X147Y121_C5Q;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_B6 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C4 = CLBLM_R_X101Y115_SLICE_X158Y115_A5Q;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C2 = CLBLM_L_X94Y121_SLICE_X148Y121_AQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C3 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C4 = CLBLM_L_X92Y120_SLICE_X145Y120_CQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C5 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_C6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C5 = CLBLL_L_X100Y118_SLICE_X157Y118_B5Q;
  assign CLBLM_R_X93Y114_SLICE_X146Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_B6 = 1'b1;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D2 = CLBLM_L_X94Y121_SLICE_X148Y121_AQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D3 = CLBLM_R_X97Y120_SLICE_X153Y120_DQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D4 = CLBLM_L_X94Y121_SLICE_X148Y121_A5Q;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D5 = CLBLM_L_X94Y121_SLICE_X148Y121_CQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_D6 = CLBLM_R_X93Y121_SLICE_X147Y121_C5Q;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B6 = CLBLM_R_X89Y117_SLICE_X140Y117_CQ;
  assign CLBLM_L_X94Y121_SLICE_X148Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C2 = CLBLM_R_X97Y131_SLICE_X152Y131_BQ;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_D1 = CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C5 = CLBLM_R_X97Y132_SLICE_X152Y132_D5Q;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_C6 = CLBLM_R_X97Y132_SLICE_X152Y132_BQ;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_D6 = CLBLM_R_X93Y129_SLICE_X147Y129_A5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A1 = CLBLM_L_X94Y113_SLICE_X148Y113_A5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A2 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A3 = CLBLM_L_X92Y113_SLICE_X144Y113_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A5 = CLBLM_R_X93Y115_SLICE_X147Y115_CO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_A6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B1 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B2 = CLBLM_L_X94Y116_SLICE_X148Y116_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B3 = CLBLM_L_X94Y115_SLICE_X148Y115_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B5 = CLBLM_R_X93Y113_SLICE_X147Y113_CO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_B6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C2 = CLBLM_L_X90Y113_SLICE_X142Y113_CO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C4 = CLBLM_L_X94Y115_SLICE_X148Y115_DO6;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C5 = CLBLM_L_X94Y114_SLICE_X149Y114_AQ;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_C6 = CLBLM_R_X97Y115_SLICE_X152Y115_A5Q;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D1 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D2 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D3 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D4 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D5 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_D6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X147Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A1 = CLBLM_R_X93Y115_SLICE_X146Y115_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A2 = CLBLM_L_X92Y113_SLICE_X145Y113_CO6;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A3 = CLBLM_R_X93Y118_SLICE_X147Y118_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A5 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_A6 = 1'b1;
  assign LIOB33_X0Y203_IOB_X0Y203_O = 1'b0;
  assign LIOB33_X0Y203_IOB_X0Y204_O = 1'b0;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B1 = CLBLM_R_X93Y118_SLICE_X147Y118_A5Q;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B3 = CLBLM_R_X93Y115_SLICE_X147Y115_B5Q;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B4 = CLBLM_L_X92Y113_SLICE_X145Y113_DO6;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B5 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_B6 = 1'b1;
  assign LIOB33_X0Y203_IOB_X0Y204_T = 1'b1;
  assign LIOB33_X0Y203_IOB_X0Y203_T = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A1 = CLBLM_L_X94Y122_SLICE_X149Y122_B5Q;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A2 = CLBLM_L_X94Y121_SLICE_X149Y121_BO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A5 = CLBLM_R_X95Y123_SLICE_X151Y123_B5Q;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_A6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C1 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C2 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B1 = CLBLM_R_X95Y123_SLICE_X150Y123_A5Q;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B3 = CLBLM_L_X94Y120_SLICE_X149Y120_A5Q;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B5 = CLBLM_L_X94Y121_SLICE_X149Y121_CO6;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_B6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D1 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D2 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D3 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D4 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D5 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_D6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C3 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_T = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_D6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_A6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_B6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_C6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D1 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D2 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D3 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D4 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D5 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X148Y122_D6 = 1'b1;
  assign LIOI3_X0Y245_OLOGIC_X0Y246_D1 = 1'b0;
  assign LIOI3_X0Y245_OLOGIC_X0Y246_T1 = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1 = 1'b1;
  assign LIOI3_X0Y245_OLOGIC_X0Y245_D1 = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = 1'b0;
  assign LIOI3_X0Y245_OLOGIC_X0Y245_T1 = 1'b1;
  assign RIOB33_X105Y51_IOB_X1Y52_O = 1'b0;
  assign RIOB33_X105Y51_IOB_X1Y51_O = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y233_OLOGIC_X0Y233_D1 = 1'b0;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = 1'b0;
  assign RIOB33_X105Y51_IOB_X1Y52_T = 1'b1;
  assign RIOB33_X105Y51_IOB_X1Y51_T = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = 1'b0;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_T1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A1 = CLBLM_L_X94Y116_SLICE_X148Y116_A5Q;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A2 = CLBLM_L_X94Y120_SLICE_X149Y120_AQ;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_A6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B3 = CLBLM_R_X93Y116_SLICE_X147Y116_AQ;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B5 = CLBLM_R_X93Y116_SLICE_X147Y116_BQ;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_B6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = 1'b0;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C1 = CLBLM_R_X93Y116_SLICE_X147Y116_BQ;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C4 = CLBLM_R_X93Y116_SLICE_X147Y116_AQ;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C5 = CLBLM_R_X93Y116_SLICE_X147Y116_B5Q;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_C6 = CLBLM_L_X94Y120_SLICE_X149Y120_AQ;
  assign LIOB33_X0Y205_IOB_X0Y205_O = 1'b0;
  assign LIOB33_X0Y205_IOB_X0Y206_O = 1'b0;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y205_IOB_X0Y206_T = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_D6 = 1'b1;
  assign LIOB33_X0Y205_IOB_X0Y205_T = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_T = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X147Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A1 = CLBLM_R_X93Y116_SLICE_X146Y116_B5Q;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A2 = CLBLM_L_X90Y115_SLICE_X143Y115_BQ;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_A6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B1 = CLBLM_R_X93Y116_SLICE_X146Y116_BQ;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B3 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B5 = CLBLM_L_X92Y115_SLICE_X145Y115_BQ;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_B6 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A1 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A2 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A3 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A4 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A5 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_A6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C5 = CLBLM_R_X93Y116_SLICE_X146Y116_B5Q;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C1 = CLBLM_L_X92Y115_SLICE_X145Y115_BQ;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B1 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B2 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B3 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B4 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B5 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_B6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D2 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C1 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D3 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C2 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D4 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C5 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C6 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D5 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C3 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_C4 = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_D6 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D1 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D2 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D3 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D4 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D5 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X149Y123_D6 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A4 = CLBLM_L_X94Y123_SLICE_X148Y123_BO6;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A5 = CLBLM_R_X95Y124_SLICE_X151Y124_DO6;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_A6 = CLBLM_L_X94Y124_SLICE_X148Y124_A5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_AX = CLBLM_L_X94Y123_SLICE_X148Y123_BO5;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B1 = CLBLM_L_X94Y123_SLICE_X148Y123_CQ;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B2 = CLBLM_L_X94Y123_SLICE_X148Y123_A5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B4 = CLBLM_L_X94Y123_SLICE_X148Y123_AQ;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B5 = CLBLM_L_X94Y123_SLICE_X148Y123_C5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_B6 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C2 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C3 = CLBLM_L_X94Y123_SLICE_X148Y123_AQ;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C4 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C5 = CLBLM_L_X94Y123_SLICE_X148Y123_CQ;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_C6 = 1'b1;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D1 = CLBLM_L_X94Y123_SLICE_X148Y123_C5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D2 = CLBLM_L_X94Y123_SLICE_X148Y123_AQ;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D3 = CLBLM_L_X92Y122_SLICE_X144Y122_C5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D4 = CLBLM_L_X94Y123_SLICE_X148Y123_A5Q;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D5 = CLBLM_L_X94Y123_SLICE_X148Y123_CQ;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y123_SLICE_X148Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y53_IOB_X1Y54_O = 1'b0;
  assign RIOB33_X105Y53_IOB_X1Y53_O = 1'b0;
  assign RIOB33_X105Y53_IOB_X1Y54_T = 1'b1;
  assign RIOB33_X105Y53_IOB_X1Y53_T = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D4 = CLBLM_R_X93Y112_SLICE_X146Y112_DO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D6 = CLBLM_R_X93Y113_SLICE_X146Y113_A5Q;
  assign LIOB33_X0Y207_IOB_X0Y208_O = 1'b0;
  assign LIOB33_X0Y207_IOB_X0Y207_O = 1'b0;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A1 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A2 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A3 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A5 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_A6 = 1'b1;
  assign LIOB33_X0Y207_IOB_X0Y207_T = 1'b1;
  assign LIOB33_X0Y207_IOB_X0Y208_T = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B1 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B2 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B3 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B5 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_B6 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C1 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C2 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C3 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A3 = CLBLM_R_X93Y113_SLICE_X146Y113_B5Q;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C5 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_C6 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D1 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D2 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D3 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D5 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X147Y117_D6 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A2 = CLBLM_R_X93Y117_SLICE_X146Y117_B5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A3 = CLBLM_R_X97Y117_SLICE_X152Y117_CO6;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A4 = CLBLM_L_X94Y116_SLICE_X149Y116_A5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A5 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_A6 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B2 = CLBLM_R_X93Y117_SLICE_X146Y117_BQ;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B3 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B5 = CLBLM_R_X93Y116_SLICE_X146Y116_AQ;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_B6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B1 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A1 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A2 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A3 = CLBLM_L_X94Y124_SLICE_X149Y124_AQ;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A5 = CLBLM_L_X98Y128_SLICE_X154Y128_AQ;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_A6 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C1 = CLBLM_R_X93Y116_SLICE_X146Y116_AQ;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B1 = CLBLM_R_X93Y124_SLICE_X147Y124_A5Q;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B3 = CLBLM_L_X92Y113_SLICE_X144Y113_AQ;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B3 = CLBLM_R_X93Y124_SLICE_X147Y124_DO6;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B5 = CLBLM_L_X94Y124_SLICE_X148Y124_AQ;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D1 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D2 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D3 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D5 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C2 = CLBLM_L_X94Y128_SLICE_X149Y128_C5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_D6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B5 = CLBLM_L_X92Y113_SLICE_X144Y113_BQ;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_B6 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C3 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C4 = CLBLM_L_X94Y124_SLICE_X149Y124_A5Q;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C6 = CLBLM_L_X98Y128_SLICE_X154Y128_AQ;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D1 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D2 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D3 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D4 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D5 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_D6 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A1 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A2 = CLBLM_L_X94Y124_SLICE_X148Y124_A5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A3 = CLBLM_R_X93Y126_SLICE_X146Y126_AQ;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A5 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_A6 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B1 = CLBLM_L_X94Y125_SLICE_X148Y125_BQ;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B3 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B4 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B5 = CLBLM_L_X94Y124_SLICE_X148Y124_BQ;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_B6 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y56_O = 1'b0;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C1 = CLBLM_L_X94Y123_SLICE_X148Y123_A5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C2 = CLBLM_L_X94Y124_SLICE_X148Y124_CQ;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C4 = CLBLM_R_X93Y125_SLICE_X147Y125_A5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C5 = CLBLM_R_X93Y124_SLICE_X146Y124_A5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_C6 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y55_O = 1'b0;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y55_IOB_X1Y56_T = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y55_T = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D2 = CLBLM_L_X94Y125_SLICE_X148Y125_BQ;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D3 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D4 = CLBLM_L_X94Y124_SLICE_X148Y124_BQ;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D5 = CLBLM_L_X94Y124_SLICE_X148Y124_B5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_D6 = CLBLM_R_X93Y124_SLICE_X147Y124_B5Q;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B2 = CLBLL_L_X100Y121_SLICE_X157Y121_C5Q;
  assign CLBLM_L_X94Y124_SLICE_X148Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B3 = CLBLL_L_X102Y121_SLICE_X160Y121_AQ;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B4 = CLBLL_L_X100Y121_SLICE_X157Y121_BQ;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B5 = CLBLL_L_X102Y120_SLICE_X160Y120_C5Q;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C3 = CLBLL_L_X102Y121_SLICE_X161Y121_DO6;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C4 = CLBLL_L_X100Y122_SLICE_X157Y122_CQ;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C6 = CLBLL_L_X102Y121_SLICE_X161Y121_C5Q;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y209_IOB_X0Y210_O = 1'b0;
  assign LIOB33_X0Y209_IOB_X0Y209_O = 1'b0;
  assign LIOI3_X0Y247_OLOGIC_X0Y248_D1 = 1'b0;
  assign LIOB33_X0Y209_IOB_X0Y210_T = 1'b1;
  assign LIOB33_X0Y209_IOB_X0Y209_T = 1'b1;
  assign LIOI3_X0Y247_OLOGIC_X0Y248_T1 = 1'b1;
  assign LIOI3_X0Y247_OLOGIC_X0Y247_D1 = 1'b0;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = 1'b0;
  assign LIOI3_X0Y247_OLOGIC_X0Y247_T1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A2 = CLBLM_L_X94Y119_SLICE_X149Y119_B5Q;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A3 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A5 = CLBLM_L_X94Y119_SLICE_X149Y119_AQ;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_A6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = 1'b0;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B2 = CLBLM_R_X93Y118_SLICE_X147Y118_BQ;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B3 = CLBLM_R_X93Y118_SLICE_X147Y118_AQ;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B5 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_B6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = 1'b0;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C1 = CLBLM_L_X94Y119_SLICE_X149Y119_AQ;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C2 = CLBLM_R_X93Y118_SLICE_X147Y118_AQ;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C3 = CLBLM_R_X93Y118_SLICE_X147Y118_BQ;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C5 = CLBLM_R_X93Y118_SLICE_X147Y118_B5Q;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_C6 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_D1 = 1'b0;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = 1'b0;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D2 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D3 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D5 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_D6 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_T1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X147Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A2 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A3 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A5 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_A6 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = 1'b0;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B2 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B3 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B5 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_B6 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A1 = CLBLM_L_X98Y126_SLICE_X155Y126_DO6;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C2 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C3 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C5 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_C6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A3 = CLBLM_L_X94Y125_SLICE_X149Y125_BO6;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A5 = CLBLM_L_X94Y127_SLICE_X149Y127_AQ;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_AX = CLBLM_L_X94Y125_SLICE_X149Y125_BO5;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B1 = CLBLM_L_X94Y125_SLICE_X149Y125_AQ;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B3 = CLBLM_L_X94Y125_SLICE_X149Y125_A5Q;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D1 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D2 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D3 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D4 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D5 = 1'b1;
  assign CLBLM_R_X93Y118_SLICE_X146Y118_D6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C4 = CLBLM_R_X95Y125_SLICE_X150Y125_BQ;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C5 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C2 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_C3 = CLBLM_L_X94Y125_SLICE_X149Y125_DQ;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D2 = CLBLM_R_X95Y128_SLICE_X150Y128_BQ;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D3 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D4 = CLBLM_L_X94Y125_SLICE_X149Y125_AQ;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D5 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_D6 = 1'b1;
  assign RIOB33_X105Y57_IOB_X1Y57_O = 1'b0;
  assign RIOB33_X105Y57_IOB_X1Y58_O = 1'b0;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A1 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A2 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A3 = CLBLM_L_X94Y125_SLICE_X148Y125_AQ;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A5 = CLBLM_L_X94Y121_SLICE_X149Y121_AQ;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_A6 = 1'b1;
  assign RIOB33_X105Y57_IOB_X1Y57_T = 1'b1;
  assign RIOB33_X105Y57_IOB_X1Y58_T = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B1 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B3 = CLBLM_L_X94Y122_SLICE_X149Y122_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B4 = CLBLM_R_X95Y126_SLICE_X150Y126_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B5 = CLBLM_L_X94Y125_SLICE_X148Y125_CO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_B6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C1 = CLBLM_R_X93Y120_SLICE_X146Y120_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C2 = CLBLM_L_X94Y125_SLICE_X148Y125_AQ;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C3 = CLBLM_R_X95Y125_SLICE_X151Y125_CO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C5 = CLBLM_L_X94Y124_SLICE_X148Y124_DO6;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D1 = CLBLM_L_X94Y125_SLICE_X149Y125_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D2 = CLBLM_L_X94Y125_SLICE_X149Y125_AQ;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D3 = CLBLM_R_X93Y125_SLICE_X147Y125_A5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D5 = CLBLM_L_X94Y125_SLICE_X149Y125_DQ;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_D6 = CLBLM_L_X94Y125_SLICE_X149Y125_C5Q;
  assign CLBLM_L_X94Y125_SLICE_X148Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C3 = CLBLM_L_X98Y113_SLICE_X154Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C5 = CLBLM_R_X93Y113_SLICE_X146Y113_DO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C6 = CLBLM_R_X97Y113_SLICE_X152Y113_BO6;
  assign LIOB33_X0Y211_IOB_X0Y212_O = 1'b0;
  assign LIOB33_X0Y211_IOB_X0Y211_O = 1'b0;
  assign LIOB33_X0Y211_IOB_X0Y212_T = 1'b1;
  assign LIOB33_X0Y211_IOB_X0Y211_T = 1'b1;
  assign LIOB33_X0Y91_IOB_X0Y92_O = 1'b0;
  assign LIOB33_X0Y91_IOB_X0Y91_O = 1'b0;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A2 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A3 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A4 = CLBLM_R_X93Y119_SLICE_X147Y119_B5Q;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A5 = CLBLM_L_X94Y122_SLICE_X149Y122_AQ;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_A6 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B2 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B3 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B4 = CLBLM_L_X94Y122_SLICE_X149Y122_BQ;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B5 = CLBLM_R_X93Y119_SLICE_X147Y119_BQ;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_B6 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C1 = CLBLM_R_X93Y119_SLICE_X147Y119_BQ;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C3 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C4 = CLBLM_R_X93Y119_SLICE_X147Y119_A5Q;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C5 = CLBLM_R_X93Y119_SLICE_X147Y119_B5Q;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_C6 = CLBLM_L_X94Y122_SLICE_X149Y122_BQ;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D1 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D2 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C4 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D3 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D4 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D5 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_D6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C5 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X147Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y91_IOB_X0Y92_T = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_C6 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A2 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A3 = CLBLM_L_X90Y119_SLICE_X143Y119_DO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A4 = CLBLM_R_X93Y119_SLICE_X146Y119_B5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A5 = CLBLM_R_X93Y119_SLICE_X146Y119_C5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_A6 = 1'b1;
  assign LIOB33_X0Y91_IOB_X0Y91_T = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B2 = CLBLM_R_X93Y114_SLICE_X146Y114_A5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B3 = CLBLM_R_X93Y119_SLICE_X147Y119_A5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B4 = CLBLM_L_X90Y118_SLICE_X143Y118_CO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B5 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_B6 = 1'b1;
  assign CLBLM_R_X93Y115_SLICE_X146Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A1 = CLBLM_L_X94Y127_SLICE_X149Y127_B5Q;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A2 = CLBLM_L_X94Y125_SLICE_X149Y125_D5Q;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A3 = CLBLM_R_X93Y125_SLICE_X147Y125_AQ;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A4 = CLBLM_L_X94Y127_SLICE_X149Y127_BQ;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C6 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_A6 = CLBLM_R_X95Y128_SLICE_X150Y128_BQ;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C1 = CLBLM_R_X93Y119_SLICE_X147Y119_AQ;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C2 = CLBLM_R_X93Y119_SLICE_X146Y119_CQ;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_B6 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D2 = CLBLM_R_X93Y119_SLICE_X146Y119_CQ;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D3 = CLBLM_R_X93Y119_SLICE_X147Y119_AQ;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_C6 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D4 = 1'b1;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D5 = CLBLM_L_X94Y122_SLICE_X149Y122_AQ;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A5 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_A6 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X149Y126_D6 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_A6 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_B6 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_C6 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D1 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D2 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D3 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D4 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D5 = 1'b1;
  assign CLBLM_L_X94Y126_SLICE_X148Y126_D6 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_B6 = CLBLM_R_X97Y132_SLICE_X152Y132_CO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C1 = CLBLM_R_X97Y132_SLICE_X152Y132_BQ;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C2 = CLBLM_R_X97Y132_SLICE_X152Y132_D5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C5 = CLBLM_R_X97Y132_SLICE_X152Y132_B5Q;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_C6 = 1'b1;
  assign LIOB33_X0Y213_IOB_X0Y214_O = 1'b0;
  assign LIOB33_X0Y213_IOB_X0Y213_O = 1'b0;
  assign LIOB33_X0Y213_IOB_X0Y214_T = 1'b1;
  assign LIOB33_X0Y213_IOB_X0Y213_T = 1'b1;
  assign CLBLM_R_X97Y132_SLICE_X152Y132_D6 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A2 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A3 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A4 = CLBLM_L_X94Y120_SLICE_X148Y120_BQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A5 = CLBLM_R_X93Y120_SLICE_X146Y120_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_A6 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B2 = CLBLM_R_X93Y120_SLICE_X147Y120_BQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B3 = CLBLM_R_X93Y120_SLICE_X147Y120_AQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B4 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B5 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_B6 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C1 = CLBLM_R_X93Y120_SLICE_X147Y120_A5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C2 = CLBLM_R_X93Y120_SLICE_X147Y120_CQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C3 = CLBLM_L_X92Y119_SLICE_X144Y119_C5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C5 = CLBLM_R_X93Y120_SLICE_X147Y120_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_C6 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D1 = CLBLM_L_X94Y120_SLICE_X148Y120_BQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D2 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D3 = CLBLM_R_X93Y120_SLICE_X147Y120_BQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D5 = CLBLM_R_X93Y120_SLICE_X147Y120_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_D6 = CLBLM_R_X93Y120_SLICE_X147Y120_AQ;
  assign CLBLM_R_X93Y120_SLICE_X147Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y61_IOB_X1Y62_O = 1'b0;
  assign RIOB33_X105Y61_IOB_X1Y61_O = 1'b0;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A2 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A3 = CLBLM_R_X93Y119_SLICE_X146Y119_A5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A4 = CLBLM_L_X92Y120_SLICE_X144Y120_CO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A5 = CLBLM_R_X93Y124_SLICE_X147Y124_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_A6 = 1'b1;
  assign RIOB33_X105Y61_IOB_X1Y61_T = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B2 = CLBLM_R_X93Y120_SLICE_X146Y120_BQ;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B3 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B4 = CLBLM_L_X94Y120_SLICE_X148Y120_CQ;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B5 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_B6 = 1'b1;
  assign RIOB33_X105Y61_IOB_X1Y62_T = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C1 = CLBLM_L_X92Y119_SLICE_X144Y119_C5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C2 = CLBLM_L_X92Y119_SLICE_X145Y119_DO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C5 = CLBLM_R_X95Y122_SLICE_X150Y122_DO6;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_C6 = CLBLM_L_X92Y120_SLICE_X144Y120_AQ;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A2 = CLBLM_L_X94Y127_SLICE_X149Y127_A5Q;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A3 = CLBLM_L_X94Y130_SLICE_X149Y130_AQ;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A4 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A5 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_A6 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B1 = CLBLM_R_X97Y126_SLICE_X153Y126_DO6;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D2 = CLBLM_R_X93Y120_SLICE_X147Y120_A5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D3 = CLBLM_R_X93Y120_SLICE_X146Y120_BQ;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D4 = 1'b1;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D5 = CLBLM_R_X93Y120_SLICE_X146Y120_B5Q;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_D6 = CLBLM_L_X94Y120_SLICE_X148Y120_CQ;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B5 = CLBLM_L_X94Y127_SLICE_X149Y127_A5Q;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_BX = CLBLM_L_X94Y127_SLICE_X149Y127_CO5;
  assign CLBLM_R_X93Y120_SLICE_X146Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C1 = CLBLM_L_X94Y125_SLICE_X149Y125_D5Q;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C2 = CLBLM_R_X95Y128_SLICE_X150Y128_BQ;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C3 = CLBLM_L_X94Y127_SLICE_X149Y127_BQ;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C5 = CLBLM_L_X94Y127_SLICE_X149Y127_B5Q;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_C6 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D1 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D2 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D4 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D5 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D6 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_D3 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = 1'b0;
  assign CLBLM_L_X94Y127_SLICE_X149Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A1 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A2 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A3 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A4 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A5 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_A6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B3 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = 1'b0;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B1 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B2 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B3 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B4 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B5 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_B6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B4 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B5 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = 1'b0;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B6 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C1 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C2 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C3 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C4 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C5 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_C6 = 1'b1;
  assign LIOI3_X0Y5_OLOGIC_X0Y6_D1 = 1'b0;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = 1'b0;
  assign LIOI3_X0Y5_OLOGIC_X0Y6_T1 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D1 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D2 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D3 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D4 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D5 = 1'b1;
  assign CLBLM_L_X94Y127_SLICE_X148Y127_D6 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_D1 = 1'b0;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign LIOI3_X0Y5_OLOGIC_X0Y5_D1 = 1'b0;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign LIOI3_X0Y5_OLOGIC_X0Y5_T1 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_D1 = 1'b0;
  assign LIOB33_X0Y215_IOB_X0Y216_O = 1'b0;
  assign LIOB33_X0Y215_IOB_X0Y215_O = 1'b0;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1 = 1'b0;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign LIOB33_X0Y215_IOB_X0Y216_T = 1'b1;
  assign LIOB33_X0Y215_IOB_X0Y215_T = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A1 = CLBLM_R_X93Y121_SLICE_X147Y121_B5Q;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A3 = CLBLM_R_X93Y121_SLICE_X147Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A4 = CLBLM_R_X93Y121_SLICE_X147Y121_AQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A5 = CLBLM_R_X93Y121_SLICE_X146Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_A6 = 1'b1;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A5 = CLBLM_R_X97Y131_SLICE_X153Y131_AQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B2 = CLBLM_L_X92Y121_SLICE_X144Y121_BQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B3 = CLBLM_R_X93Y121_SLICE_X147Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B4 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B5 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_B6 = 1'b1;
  assign RIOB33_X105Y63_IOB_X1Y63_O = 1'b0;
  assign RIOB33_X105Y63_IOB_X1Y64_O = 1'b0;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C1 = CLBLM_R_X93Y121_SLICE_X146Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C2 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C3 = CLBLM_L_X94Y121_SLICE_X148Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C5 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_C6 = 1'b1;
  assign RIOB33_X105Y63_IOB_X1Y64_T = 1'b1;
  assign RIOB33_X105Y63_IOB_X1Y63_T = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y131_SLICE_X152Y131_A6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D1 = CLBLM_R_X97Y120_SLICE_X153Y120_D5Q;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D2 = CLBLM_R_X93Y121_SLICE_X147Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D4 = CLBLM_R_X93Y121_SLICE_X146Y121_CQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D5 = CLBLM_R_X93Y121_SLICE_X147Y121_B5Q;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_D6 = CLBLM_R_X93Y121_SLICE_X147Y121_AQ;
  assign CLBLM_R_X93Y121_SLICE_X147Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A2 = CLBLM_R_X93Y121_SLICE_X146Y121_A5Q;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A3 = CLBLM_L_X92Y119_SLICE_X145Y119_AQ;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A4 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A5 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_A6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B2 = CLBLM_R_X93Y121_SLICE_X146Y121_BQ;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B3 = CLBLM_R_X93Y122_SLICE_X147Y122_C5Q;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B4 = CLBLM_R_X93Y121_SLICE_X147Y121_BQ;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B5 = CLBLM_L_X92Y121_SLICE_X144Y121_BQ;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_B6 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A1 = CLBLM_R_X97Y128_SLICE_X153Y128_DO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A4 = CLBLM_L_X94Y128_SLICE_X149Y128_BO6;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A5 = CLBLM_L_X94Y130_SLICE_X149Y130_AQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C1 = CLBLM_R_X93Y121_SLICE_X146Y121_A5Q;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C2 = CLBLM_R_X93Y121_SLICE_X147Y121_AO6;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_AX = CLBLM_L_X94Y128_SLICE_X149Y128_BO5;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B2 = CLBLM_L_X94Y128_SLICE_X149Y128_A5Q;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B3 = CLBLM_L_X94Y128_SLICE_X149Y128_AQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B4 = CLBLM_L_X94Y128_SLICE_X149Y128_CQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B5 = CLBLM_L_X94Y129_SLICE_X148Y129_B5Q;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_B6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D2 = CLBLM_R_X93Y122_SLICE_X147Y122_C5Q;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D3 = CLBLM_R_X93Y121_SLICE_X146Y121_BQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C1 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D5 = CLBLM_R_X97Y121_SLICE_X153Y121_CQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C3 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D6 = CLBLM_R_X93Y121_SLICE_X147Y121_BQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C4 = CLBLM_L_X94Y124_SLICE_X149Y124_A5Q;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C5 = CLBLM_L_X94Y128_SLICE_X149Y128_AQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_C6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D2 = CLBLM_R_X93Y128_SLICE_X147Y128_DQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D3 = CLBLM_L_X94Y129_SLICE_X148Y129_B5Q;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D4 = CLBLM_L_X94Y128_SLICE_X149Y128_A5Q;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D5 = CLBLM_L_X94Y128_SLICE_X149Y128_AQ;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_D6 = CLBLM_L_X94Y128_SLICE_X149Y128_CQ;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C3 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X149Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C4 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A1 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A2 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A3 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A4 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A5 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_A6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C5 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C6 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B1 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B2 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B3 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B4 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B5 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_B6 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C1 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C2 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C3 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C4 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C5 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_C6 = 1'b1;
  assign LIOB33_X0Y217_IOB_X0Y218_O = 1'b0;
  assign LIOB33_X0Y217_IOB_X0Y217_O = 1'b0;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D1 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D2 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D3 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D4 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D5 = 1'b1;
  assign CLBLM_L_X94Y128_SLICE_X148Y128_D6 = 1'b1;
  assign LIOB33_X0Y217_IOB_X0Y218_T = 1'b1;
  assign LIOB33_X0Y217_IOB_X0Y217_T = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D2 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = 1'b0;
  assign RIOB33_X105Y65_IOB_X1Y66_O = 1'b0;
  assign RIOB33_X105Y65_IOB_X1Y65_O = 1'b0;
  assign RIOB33_X105Y65_IOB_X1Y66_T = 1'b1;
  assign RIOB33_X105Y65_IOB_X1Y65_T = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A1 = CLBLM_L_X92Y121_SLICE_X144Y121_AQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A4 = CLBLM_R_X93Y122_SLICE_X147Y122_BO6;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_A6 = CLBLM_L_X90Y124_SLICE_X142Y124_DO6;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_AX = CLBLM_R_X93Y122_SLICE_X147Y122_BO5;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B1 = CLBLM_R_X93Y122_SLICE_X147Y122_AQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B2 = CLBLM_R_X93Y123_SLICE_X147Y123_C5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B4 = CLBLM_R_X93Y122_SLICE_X147Y122_CQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B5 = CLBLM_R_X93Y122_SLICE_X147Y122_A5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_B6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C2 = CLBLM_R_X93Y121_SLICE_X147Y121_BQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C3 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C5 = CLBLM_R_X93Y122_SLICE_X147Y122_AQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_C6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D2 = CLBLM_R_X93Y123_SLICE_X147Y123_C5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D3 = CLBLM_R_X97Y121_SLICE_X153Y121_C5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D4 = CLBLM_R_X93Y122_SLICE_X147Y122_A5Q;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D5 = CLBLM_R_X93Y122_SLICE_X147Y122_AQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_D6 = CLBLM_R_X93Y122_SLICE_X147Y122_CQ;
  assign CLBLM_R_X93Y122_SLICE_X147Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A1 = CLBLM_L_X92Y123_SLICE_X145Y123_BQ;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A3 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A4 = CLBLM_R_X93Y123_SLICE_X146Y123_BQ;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_A6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B1 = CLBLM_L_X92Y123_SLICE_X145Y123_BQ;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B2 = CLBLM_R_X97Y123_SLICE_X152Y123_C5Q;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B3 = CLBLM_R_X93Y122_SLICE_X146Y122_AQ;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B4 = CLBLM_L_X92Y122_SLICE_X145Y122_B5Q;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_B6 = CLBLM_L_X92Y122_SLICE_X145Y122_AQ;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A1 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C3 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C4 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C5 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C6 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A3 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A5 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_A6 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B1 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B2 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B3 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_B4 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D3 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C1 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C2 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D5 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C3 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_D6 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C5 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_C6 = 1'b1;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B3 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D1 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D2 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D3 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D5 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X149Y129_D6 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A1 = CLBLM_L_X94Y129_SLICE_X148Y129_AQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A2 = CLBLM_L_X94Y129_SLICE_X148Y129_BQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A4 = CLBLM_R_X95Y129_SLICE_X150Y129_C5Q;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A5 = CLBLM_L_X94Y130_SLICE_X148Y130_AQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_A6 = 1'b1;
  assign LIOB33_X0Y219_IOB_X0Y219_O = 1'b0;
  assign LIOB33_X0Y219_IOB_X0Y220_O = 1'b0;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B1 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B2 = CLBLM_L_X94Y128_SLICE_X149Y128_CQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B5 = CLBLM_L_X94Y130_SLICE_X148Y130_AQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_B6 = 1'b1;
  assign LIOB33_X0Y219_IOB_X0Y219_T = 1'b1;
  assign LIOB33_X0Y219_IOB_X0Y220_T = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C1 = CLBLM_R_X101Y110_SLICE_X158Y110_BQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C1 = CLBLM_L_X94Y130_SLICE_X148Y130_AQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C2 = CLBLM_L_X94Y129_SLICE_X148Y129_AQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C3 = CLBLM_R_X95Y129_SLICE_X150Y129_C5Q;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C5 = CLBLM_L_X94Y129_SLICE_X148Y129_BQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_C6 = CLBLM_R_X93Y128_SLICE_X147Y128_A5Q;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C2 = CLBLL_L_X100Y111_SLICE_X157Y111_CQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B2 = CLBLL_L_X102Y122_SLICE_X160Y122_B5Q;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B3 = CLBLL_L_X102Y124_SLICE_X160Y124_AQ;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D1 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D2 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D3 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D4 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D5 = 1'b1;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_D6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B4 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C4 = CLBLM_R_X101Y110_SLICE_X158Y110_A5Q;
  assign CLBLM_L_X94Y129_SLICE_X148Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C1 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C2 = CLBLL_L_X102Y122_SLICE_X161Y122_A5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_TBYTETERM_X0Y237_OLOGIC_X0Y238_D1 = 1'b0;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C4 = CLBLL_L_X102Y123_SLICE_X161Y123_A5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C5 = CLBLM_R_X101Y122_SLICE_X158Y122_CO6;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_C6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = 1'b0;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = 1'b0;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = 1'b0;
  assign RIOB33_X105Y67_IOB_X1Y68_O = 1'b0;
  assign RIOB33_X105Y67_IOB_X1Y67_O = 1'b0;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_D1 = 1'b0;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign RIOB33_X105Y67_IOB_X1Y68_T = 1'b1;
  assign RIOB33_X105Y67_IOB_X1Y67_T = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_T1 = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1 = 1'b0;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A1 = CLBLM_R_X93Y123_SLICE_X147Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A2 = CLBLM_R_X93Y123_SLICE_X146Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A4 = CLBLM_R_X93Y123_SLICE_X147Y123_B5Q;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A5 = CLBLM_L_X92Y123_SLICE_X144Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_A6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B1 = CLBLM_R_X93Y123_SLICE_X147Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B3 = CLBLM_L_X92Y123_SLICE_X144Y123_BQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B4 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B5 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1 = 1'b0;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C1 = CLBLM_L_X92Y123_SLICE_X144Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C3 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C4 = CLBLM_R_X93Y122_SLICE_X147Y122_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C5 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D1 = CLBLM_L_X92Y123_SLICE_X144Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D2 = CLBLM_R_X93Y123_SLICE_X147Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D4 = CLBLM_R_X93Y123_SLICE_X146Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D5 = CLBLM_R_X93Y123_SLICE_X147Y123_B5Q;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_D6 = CLBLM_R_X97Y123_SLICE_X153Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X147Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A1 = CLBLM_R_X93Y123_SLICE_X146Y123_B5Q;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A2 = CLBLM_R_X93Y123_SLICE_X146Y123_AQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A3 = CLBLM_R_X93Y123_SLICE_X147Y123_BQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A5 = CLBLM_L_X92Y123_SLICE_X144Y123_BQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_A6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B1 = CLBLM_L_X92Y123_SLICE_X145Y123_CQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B2 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B3 = CLBLM_R_X93Y123_SLICE_X147Y123_BQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B5 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_B6 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A1 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A2 = CLBLM_R_X95Y132_SLICE_X151Y132_AQ;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A4 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A5 = CLBLM_L_X94Y130_SLICE_X149Y130_A5Q;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_A6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C6 = CLBLM_L_X92Y123_SLICE_X145Y123_B5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D2 = CLBLM_L_X98Y131_SLICE_X154Y131_CQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D3 = CLBLM_L_X98Y131_SLICE_X154Y131_AQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B1 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B2 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B3 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B5 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_B6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_CX = CLBLM_R_X93Y123_SLICE_X147Y123_AO5;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D1 = CLBLM_L_X92Y123_SLICE_X144Y123_BQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D2 = CLBLM_R_X93Y123_SLICE_X146Y123_AQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D3 = CLBLM_R_X97Y123_SLICE_X153Y123_C5Q;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C1 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C2 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D5 = CLBLM_R_X93Y123_SLICE_X146Y123_B5Q;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C3 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_D6 = CLBLM_R_X93Y123_SLICE_X147Y123_BQ;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C4 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C5 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_C6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y221_IOB_X0Y221_T = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D1 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D2 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D3 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D4 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D5 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_D6 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X149Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A1 = CLBLM_R_X95Y131_SLICE_X150Y131_A5Q;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A2 = CLBLM_L_X94Y129_SLICE_X148Y129_AO6;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_A6 = CLBLM_R_X97Y130_SLICE_X152Y130_CO6;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B1 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B2 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B3 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B4 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B5 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_B6 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C1 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C2 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C3 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C4 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C5 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_C6 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D1 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D2 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D3 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D4 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D5 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_D6 = 1'b1;
  assign CLBLM_L_X94Y130_SLICE_X148Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C4 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C5 = CLBLM_R_X95Y115_SLICE_X150Y115_B5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y69_IOB_X1Y70_O = 1'b0;
  assign RIOB33_X105Y69_IOB_X1Y69_O = 1'b0;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A5 = CLBLM_R_X101Y131_SLICE_X158Y131_CO6;
  assign RIOB33_X105Y69_IOB_X1Y70_T = 1'b1;
  assign RIOB33_X105Y69_IOB_X1Y69_T = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_D1 = 1'b0;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B4 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B5 = CLBLM_R_X101Y131_SLICE_X159Y131_AQ;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B6 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A1 = CLBLM_R_X93Y120_SLICE_X146Y120_CO6;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A3 = CLBLM_R_X93Y120_SLICE_X146Y120_A5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A4 = CLBLM_L_X94Y124_SLICE_X148Y124_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A5 = CLBLM_R_X93Y124_SLICE_X147Y124_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_A6 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B1 = CLBLM_R_X95Y124_SLICE_X150Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B3 = CLBLM_L_X94Y124_SLICE_X148Y124_B5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B4 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B5 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_B6 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A5 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A6 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C1 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C3 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C4 = CLBLM_R_X93Y124_SLICE_X147Y124_BQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C5 = CLBLM_R_X93Y124_SLICE_X147Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_C6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C1 = CLBLM_R_X101Y131_SLICE_X159Y131_AQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D1 = CLBLM_R_X93Y124_SLICE_X147Y124_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D2 = CLBLM_R_X93Y124_SLICE_X147Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D3 = CLBLM_R_X93Y124_SLICE_X147Y124_BQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D4 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D5 = CLBLM_R_X95Y124_SLICE_X150Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C3 = CLBLM_R_X93Y116_SLICE_X146Y116_BQ;
  assign CLBLM_R_X93Y124_SLICE_X147Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B2 = CLBLL_L_X100Y120_SLICE_X157Y120_BQ;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C4 = CLBLM_R_X93Y116_SLICE_X146Y116_A5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A1 = CLBLM_R_X95Y125_SLICE_X150Y125_DO6;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A2 = CLBLM_R_X93Y126_SLICE_X146Y126_AQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A4 = CLBLM_R_X93Y124_SLICE_X146Y124_BO6;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B4 = CLBLL_L_X100Y119_SLICE_X156Y119_BQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_AX = CLBLM_R_X93Y124_SLICE_X146Y124_BO5;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_C6 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B1 = CLBLM_R_X93Y124_SLICE_X146Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B2 = CLBLM_R_X93Y124_SLICE_X146Y124_A5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B3 = CLBLM_R_X93Y124_SLICE_X146Y124_AQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B5 = CLBLM_R_X93Y124_SLICE_X146Y124_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_B6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X153Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y223_IOB_X0Y223_O = 1'b0;
  assign LIOB33_X0Y223_IOB_X0Y224_O = 1'b0;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C1 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C2 = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C3 = CLBLM_R_X93Y124_SLICE_X146Y124_AQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C5 = CLBLM_R_X93Y124_SLICE_X146Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_C6 = 1'b1;
  assign LIOB33_X0Y223_IOB_X0Y223_T = 1'b1;
  assign CLBLM_R_X93Y116_SLICE_X146Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y223_IOB_X0Y224_T = 1'b1;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D1 = CLBLM_R_X93Y124_SLICE_X146Y124_C5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D2 = CLBLM_R_X93Y124_SLICE_X146Y124_AQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D3 = CLBLM_L_X92Y122_SLICE_X144Y122_CQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D4 = CLBLM_R_X93Y124_SLICE_X146Y124_A5Q;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D5 = CLBLM_R_X93Y124_SLICE_X146Y124_CQ;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y124_SLICE_X146Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A1 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A2 = CLBLM_R_X89Y118_SLICE_X140Y118_A5Q;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOB33_X0Y237_IOB_X0Y238_O = 1'b0;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y237_IOB_X0Y237_O = 1'b0;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_B6 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B4 = CLBLL_R_X87Y118_SLICE_X139Y118_BO6;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOB33_X0Y237_IOB_X0Y238_T = 1'b1;
  assign LIOB33_X0Y237_IOB_X0Y237_T = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C1 = 1'b1;
  assign LIOI3_X0Y211_OLOGIC_X0Y211_D1 = 1'b0;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C2 = 1'b1;
  assign RIOB33_X105Y71_IOB_X1Y72_O = 1'b0;
  assign RIOB33_X105Y71_IOB_X1Y71_O = 1'b0;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C5 = CLBLM_R_X97Y133_SLICE_X152Y133_CQ;
  assign RIOB33_X105Y71_IOB_X1Y72_T = 1'b1;
  assign RIOB33_X105Y71_IOB_X1Y71_T = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_C6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_D6 = CLBLM_R_X97Y133_SLICE_X152Y133_AQ;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A1 = CLBLM_R_X93Y125_SLICE_X146Y125_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A3 = CLBLM_R_X93Y125_SLICE_X147Y125_AQ;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A4 = CLBLM_L_X92Y125_SLICE_X145Y125_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A5 = CLBLM_R_X93Y128_SLICE_X147Y128_DQ;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_A6 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B1 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B2 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B3 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B4 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B5 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_B6 = 1'b1;
  assign CLBLM_R_X97Y133_SLICE_X152Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C1 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C2 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C3 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C4 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C5 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign LIOB33_X0Y225_IOB_X0Y226_O = 1'b0;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y225_IOB_X0Y225_O = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D1 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D2 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D3 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D4 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D5 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_D6 = 1'b1;
  assign LIOB33_X0Y225_IOB_X0Y225_T = 1'b1;
  assign LIOB33_X0Y225_IOB_X0Y226_T = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X147Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = 1'b0;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A1 = CLBLM_R_X93Y126_SLICE_X146Y126_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A3 = CLBLM_L_X94Y125_SLICE_X148Y125_DO6;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A4 = CLBLM_R_X93Y125_SLICE_X146Y125_BO6;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_AX = CLBLM_R_X93Y125_SLICE_X146Y125_BO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B1 = CLBLM_R_X93Y125_SLICE_X146Y125_CQ;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B2 = CLBLM_R_X93Y125_SLICE_X146Y125_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B3 = CLBLM_R_X93Y125_SLICE_X146Y125_AQ;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B5 = CLBLM_R_X93Y125_SLICE_X146Y125_C5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_B6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = 1'b0;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A1 = CLBLM_R_X95Y132_SLICE_X151Y132_CQ;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A2 = CLBLM_R_X95Y132_SLICE_X150Y132_C5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A3 = CLBLM_R_X97Y132_SLICE_X152Y132_DQ;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A5 = CLBLM_R_X95Y132_SLICE_X151Y132_B5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C5 = CLBLM_R_X93Y125_SLICE_X146Y125_CQ;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C6 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_A6 = CLBLM_R_X93Y131_SLICE_X147Y131_A5Q;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B3 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B4 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_B6 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D2 = CLBLM_R_X93Y125_SLICE_X146Y125_CQ;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D3 = CLBLM_R_X93Y125_SLICE_X146Y125_AQ;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D4 = CLBLM_R_X93Y125_SLICE_X146Y125_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C3 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C4 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D6 = CLBLM_L_X90Y124_SLICE_X143Y124_C5Q;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_C6 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1 = CLBLM_R_X101Y120_SLICE_X159Y120_CO6;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D3 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D4 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X149Y132_D6 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A3 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A4 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_A6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1 = CLBLL_L_X102Y119_SLICE_X161Y119_CO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B2 = CLBLM_R_X95Y111_SLICE_X150Y111_AQ;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B4 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B6 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_B3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C3 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C4 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_C6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D1 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D2 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D3 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D4 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D5 = 1'b1;
  assign CLBLM_L_X94Y132_SLICE_X148Y132_D6 = 1'b1;
  assign RIOB33_X105Y73_IOB_X1Y74_O = 1'b0;
  assign RIOB33_X105Y73_IOB_X1Y73_O = 1'b0;
  assign RIOB33_X105Y73_IOB_X1Y74_T = 1'b1;
  assign RIOB33_X105Y73_IOB_X1Y73_T = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C4 = CLBLM_L_X98Y111_SLICE_X155Y111_BQ;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C5 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C6 = 1'b1;
  assign LIOB33_X0Y227_IOB_X0Y228_O = 1'b0;
  assign LIOB33_X0Y227_IOB_X0Y227_O = 1'b0;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A1 = CLBLM_R_X95Y129_SLICE_X150Y129_DO6;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A2 = CLBLM_L_X94Y125_SLICE_X148Y125_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A4 = CLBLM_R_X93Y126_SLICE_X147Y126_BO6;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_AX = CLBLM_R_X93Y126_SLICE_X147Y126_BO5;
  assign LIOB33_X0Y227_IOB_X0Y227_T = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B1 = CLBLM_R_X93Y126_SLICE_X147Y126_CQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B2 = CLBLM_R_X93Y126_SLICE_X147Y126_C5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B3 = CLBLM_R_X93Y126_SLICE_X147Y126_AQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B4 = CLBLM_R_X93Y126_SLICE_X147Y126_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_B6 = 1'b1;
  assign LIOB33_X0Y227_IOB_X0Y228_T = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C2 = CLBLM_R_X93Y126_SLICE_X147Y126_CQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C3 = CLBLM_R_X93Y126_SLICE_X147Y126_AQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C4 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C5 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_C6 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D1 = CLBLM_R_X93Y126_SLICE_X147Y126_C5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D2 = CLBLM_R_X93Y126_SLICE_X147Y126_CQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D4 = CLBLM_R_X93Y126_SLICE_X147Y126_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D5 = CLBLM_R_X93Y126_SLICE_X147Y126_AQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_D6 = CLBLM_L_X90Y125_SLICE_X143Y125_BQ;
  assign CLBLM_R_X93Y126_SLICE_X147Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A1 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A3 = CLBLM_R_X93Y127_SLICE_X146Y127_AQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A4 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A5 = CLBLM_R_X93Y126_SLICE_X146Y126_A5Q;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_A6 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B1 = CLBLM_R_X93Y126_SLICE_X146Y126_CQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B2 = CLBLM_R_X93Y126_SLICE_X146Y126_BQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B4 = CLBLM_R_X93Y129_SLICE_X146Y129_CQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B5 = CLBLM_R_X93Y126_SLICE_X146Y126_C5Q;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_B6 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C1 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C2 = CLBLM_R_X93Y126_SLICE_X146Y126_CQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C3 = CLBLM_R_X93Y129_SLICE_X146Y129_CQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C5 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_C6 = 1'b1;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D1 = CLBLM_R_X93Y126_SLICE_X146Y126_C5Q;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D2 = CLBLM_R_X93Y126_SLICE_X146Y126_CQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D3 = CLBLM_R_X93Y126_SLICE_X146Y126_BQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D4 = CLBLM_R_X93Y129_SLICE_X146Y129_CQ;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_D6 = CLBLM_L_X92Y126_SLICE_X145Y126_C5Q;
  assign CLBLM_R_X93Y126_SLICE_X146Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A1 = CLBLM_L_X90Y113_SLICE_X143Y113_B5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A2 = CLBLM_L_X90Y113_SLICE_X142Y113_BO6;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A3 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A5 = CLBLM_L_X92Y113_SLICE_X145Y113_A5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_A6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C2 = CLBLM_L_X98Y111_SLICE_X154Y111_AQ;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B1 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B2 = CLBLM_R_X93Y114_SLICE_X146Y114_AQ;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B3 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B5 = CLBLM_L_X90Y113_SLICE_X143Y113_C5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_B6 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C5 = CLBLM_L_X98Y111_SLICE_X154Y111_B5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C2 = CLBLM_L_X90Y113_SLICE_X143Y113_CQ;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C3 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C4 = CLBLM_R_X93Y114_SLICE_X146Y114_BQ;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C5 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_C6 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y75_IOB_X1Y76_O = 1'b0;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D1 = CLBLM_L_X90Y113_SLICE_X143Y113_C5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D2 = CLBLM_L_X90Y113_SLICE_X143Y113_CQ;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D3 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D5 = CLBLM_L_X90Y113_SLICE_X143Y113_B5Q;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_D6 = CLBLM_R_X93Y114_SLICE_X146Y114_BQ;
  assign RIOB33_X105Y75_IOB_X1Y75_O = 1'b0;
  assign CLBLM_L_X90Y113_SLICE_X143Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y75_IOB_X1Y75_T = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A1 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A3 = CLBLM_L_X90Y113_SLICE_X142Y113_AQ;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A4 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A5 = CLBLM_L_X90Y113_SLICE_X143Y113_AQ;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_A6 = 1'b1;
  assign RIOB33_X105Y75_IOB_X1Y76_T = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B2 = CLBLM_L_X92Y114_SLICE_X144Y114_DO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B4 = CLBLM_L_X90Y114_SLICE_X142Y114_B5Q;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B5 = CLBLM_L_X92Y115_SLICE_X145Y115_B5Q;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_B6 = CLBLM_L_X90Y113_SLICE_X142Y113_CO6;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C1 = CLBLM_L_X90Y113_SLICE_X143Y113_AQ;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C2 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C3 = CLBLM_L_X90Y113_SLICE_X142Y113_AQ;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C4 = CLBLM_L_X90Y113_SLICE_X142Y113_A5Q;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C5 = CLBLM_L_X90Y114_SLICE_X143Y114_A5Q;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = 1'b0;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D1 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D2 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D3 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D4 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D5 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_D6 = 1'b1;
  assign CLBLM_L_X90Y113_SLICE_X142Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C4 = CLBLM_R_X93Y117_SLICE_X146Y117_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C5 = CLBLM_L_X92Y115_SLICE_X145Y115_AQ;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C6 = CLBLM_R_X93Y117_SLICE_X146Y117_CO6;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_D1 = CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  assign LIOB33_X0Y229_IOB_X0Y230_O = 1'b0;
  assign LIOB33_X0Y229_IOB_X0Y229_O = 1'b0;
  assign LIOB33_X0Y229_IOB_X0Y230_T = 1'b1;
  assign LIOB33_X0Y229_IOB_X0Y229_T = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A2 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A3 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A4 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A5 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_A6 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B2 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B3 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B4 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B5 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_B6 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C2 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C3 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C4 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C5 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_C6 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D2 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D3 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D4 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D5 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X147Y127_D6 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A2 = CLBLM_R_X93Y127_SLICE_X146Y127_A5Q;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A3 = CLBLM_R_X93Y130_SLICE_X146Y130_AQ;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A5 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_A6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A6 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B4 = CLBLM_L_X92Y127_SLICE_X145Y127_AO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B5 = CLBLM_R_X93Y130_SLICE_X146Y130_AQ;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_B6 = CLBLM_R_X95Y128_SLICE_X150Y128_CO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C2 = CLBLM_R_X93Y129_SLICE_X146Y129_B5Q;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C3 = CLBLM_L_X92Y126_SLICE_X145Y126_AO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C4 = CLBLM_R_X95Y128_SLICE_X151Y128_AO6;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_O = 1'b0;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_T = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D1 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D2 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D3 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D4 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D5 = 1'b1;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_D6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B1 = CLBLM_R_X101Y111_SLICE_X158Y111_BQ;
  assign CLBLM_R_X93Y127_SLICE_X146Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B3 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B4 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A1 = CLBLM_L_X90Y113_SLICE_X142Y113_A5Q;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A2 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A4 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A5 = CLBLM_L_X92Y114_SLICE_X144Y114_AQ;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_A6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B5 = CLBLM_R_X101Y110_SLICE_X158Y110_AQ;
  assign RIOB33_X105Y77_IOB_X1Y77_O = 1'b0;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B1 = CLBLM_L_X90Y114_SLICE_X143Y114_AQ;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B2 = CLBLM_L_X90Y114_SLICE_X143Y114_BQ;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B4 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B5 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_B6 = 1'b1;
  assign RIOB33_X105Y77_IOB_X1Y77_T = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C1 = CLBLM_L_X90Y118_SLICE_X143Y118_DO6;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C4 = CLBLM_L_X90Y115_SLICE_X143Y115_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C5 = CLBLM_L_X90Y114_SLICE_X143Y114_DO6;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_C6 = CLBLM_L_X90Y114_SLICE_X142Y114_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = 1'b0;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D1 = CLBLM_L_X90Y114_SLICE_X143Y114_BQ;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D2 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D4 = CLBLM_L_X90Y114_SLICE_X143Y114_AQ;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D5 = CLBLM_L_X90Y114_SLICE_X143Y114_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_D6 = CLBLM_L_X92Y114_SLICE_X144Y114_AQ;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X143Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C2 = CLBLM_R_X101Y110_SLICE_X158Y110_CO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = 1'b0;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A1 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A2 = CLBLM_L_X90Y114_SLICE_X142Y114_BQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A3 = CLBLM_L_X90Y114_SLICE_X142Y114_AQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A4 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_A6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C3 = CLBLM_L_X98Y111_SLICE_X154Y111_CO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C4 = CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = 1'b0;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B1 = CLBLM_L_X90Y114_SLICE_X142Y114_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B2 = CLBLM_R_X93Y112_SLICE_X147Y112_AQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B3 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B4 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_B6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = 1'b0;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C2 = CLBLM_L_X90Y114_SLICE_X142Y114_CQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C3 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C4 = CLBLM_L_X90Y115_SLICE_X143Y115_CQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C5 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_C6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_D1 = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C4 = CLBLL_L_X102Y124_SLICE_X160Y124_CQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D1 = CLBLM_L_X90Y114_SLICE_X142Y114_C5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D2 = CLBLM_L_X90Y114_SLICE_X142Y114_CQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D3 = CLBLM_R_X89Y114_SLICE_X141Y114_A5Q;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C5 = CLBLL_L_X102Y123_SLICE_X160Y123_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D4 = CLBLM_L_X90Y115_SLICE_X143Y115_CQ;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_D6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_T1 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C6 = CLBLL_L_X102Y122_SLICE_X160Y122_B5Q;
  assign CLBLM_L_X90Y114_SLICE_X142Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1 = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_T1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1 = CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D5 = CLBLM_R_X101Y111_SLICE_X158Y111_B5Q;
  assign LIOB33_X0Y231_IOB_X0Y232_O = 1'b0;
  assign LIOB33_X0Y231_IOB_X0Y231_O = 1'b0;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D1 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D2 = CLBLL_L_X102Y123_SLICE_X160Y123_AQ;
  assign LIOB33_X0Y231_IOB_X0Y232_T = 1'b1;
  assign LIOB33_X0Y231_IOB_X0Y231_T = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D3 = CLBLL_L_X102Y123_SLICE_X160Y123_BQ;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D4 = CLBLL_L_X102Y124_SLICE_X160Y124_CQ;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D5 = CLBLL_L_X102Y123_SLICE_X160Y123_B5Q;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C2 = CLBLM_L_X98Y132_SLICE_X154Y132_CQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A1 = CLBLM_R_X93Y120_SLICE_X146Y120_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A2 = CLBLM_R_X93Y126_SLICE_X147Y126_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A4 = CLBLM_L_X92Y128_SLICE_X145Y128_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C3 = CLBLM_L_X98Y132_SLICE_X154Y132_AQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A5 = CLBLM_R_X93Y129_SLICE_X147Y129_AQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_A6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B1 = CLBLM_L_X92Y126_SLICE_X144Y126_AQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B2 = CLBLM_R_X93Y128_SLICE_X147Y128_BQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B4 = CLBLM_R_X93Y128_SLICE_X147Y128_AQ;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C5 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B5 = CLBLM_R_X93Y126_SLICE_X146Y126_BQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_B6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C6 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C1 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C3 = CLBLM_L_X92Y127_SLICE_X145Y127_AQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C4 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C5 = CLBLM_R_X93Y131_SLICE_X147Y131_B5Q;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_C6 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D1 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D3 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D4 = CLBLM_R_X93Y120_SLICE_X146Y120_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D5 = CLBLM_R_X93Y128_SLICE_X147Y128_CQ;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_D6 = CLBLM_R_X93Y128_SLICE_X146Y128_A5Q;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X147Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C2 = CLBLL_L_X100Y121_SLICE_X156Y121_CQ;
  assign LIOB33_SING_X0Y50_IOB_X0Y50_O = 1'b0;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A1 = CLBLM_L_X94Y128_SLICE_X149Y128_DO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A4 = CLBLM_R_X93Y128_SLICE_X146Y128_BO6;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A5 = CLBLM_R_X93Y127_SLICE_X146Y127_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C4 = CLBLM_R_X101Y121_SLICE_X159Y121_B5Q;
  assign LIOB33_SING_X0Y50_IOB_X0Y50_T = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_AX = CLBLM_R_X93Y128_SLICE_X146Y128_BO5;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C5 = CLBLM_R_X97Y121_SLICE_X152Y121_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B1 = CLBLM_R_X93Y128_SLICE_X146Y128_CQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B2 = CLBLM_R_X93Y128_SLICE_X146Y128_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B4 = CLBLM_R_X93Y128_SLICE_X146Y128_AQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B5 = CLBLM_R_X93Y128_SLICE_X146Y128_C5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_B6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C6 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C2 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C3 = CLBLM_R_X93Y128_SLICE_X146Y128_AQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C4 = 1'b1;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C5 = CLBLM_R_X93Y128_SLICE_X146Y128_CQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_C6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D1 = CLBLM_L_X98Y132_SLICE_X154Y132_C5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOB33_X105Y79_IOB_X1Y80_O = CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  assign RIOB33_X105Y79_IOB_X1Y79_O = 1'b0;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D3 = CLBLM_L_X98Y132_SLICE_X154Y132_AQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D1 = CLBLM_R_X93Y128_SLICE_X146Y128_C5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D2 = CLBLM_R_X93Y128_SLICE_X146Y128_CQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D3 = CLBLM_R_X93Y128_SLICE_X146Y128_AQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D4 = CLBLM_R_X93Y128_SLICE_X146Y128_A5Q;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D5 = CLBLM_L_X90Y125_SLICE_X143Y125_DQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D4 = CLBLM_L_X98Y132_SLICE_X154Y132_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D5 = CLBLM_R_X97Y132_SLICE_X153Y132_CQ;
  assign CLBLM_R_X93Y128_SLICE_X146Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y79_IOB_X1Y79_T = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D6 = CLBLM_L_X98Y132_SLICE_X154Y132_CQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D4 = CLBLM_L_X90Y117_SLICE_X142Y117_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A1 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A2 = CLBLM_R_X89Y117_SLICE_X140Y117_AQ;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A4 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A5 = CLBLM_L_X90Y115_SLICE_X143Y115_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_A6 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B1 = CLBLM_L_X92Y115_SLICE_X145Y115_CO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B2 = CLBLM_L_X90Y114_SLICE_X143Y114_B5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B4 = CLBLM_L_X92Y115_SLICE_X145Y115_B5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B5 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_B6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C2 = CLBLM_L_X90Y115_SLICE_X142Y115_CO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C3 = CLBLM_L_X92Y114_SLICE_X144Y114_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C4 = CLBLM_L_X90Y117_SLICE_X143Y117_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C5 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_C6 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A1 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A2 = CLBLL_L_X100Y111_SLICE_X156Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A3 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A5 = CLBLL_L_X100Y111_SLICE_X157Y111_AQ;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D1 = CLBLM_R_X89Y115_SLICE_X141Y115_DO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D2 = CLBLM_R_X89Y114_SLICE_X141Y114_CO6;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D4 = CLBLM_L_X90Y115_SLICE_X143Y115_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_D6 = CLBLM_R_X89Y115_SLICE_X141Y115_CQ;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B1 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X143Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B2 = CLBLL_L_X100Y111_SLICE_X156Y111_BQ;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B3 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A1 = CLBLM_L_X90Y115_SLICE_X143Y115_B5Q;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A2 = CLBLM_L_X90Y115_SLICE_X143Y115_DO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A4 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A5 = CLBLM_R_X89Y114_SLICE_X141Y114_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_A6 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C2 = CLBLM_R_X101Y111_SLICE_X159Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B2 = CLBLM_L_X90Y116_SLICE_X142Y116_BO6;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B4 = CLBLM_R_X89Y117_SLICE_X140Y117_AQ;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_B6 = CLBLM_R_X89Y115_SLICE_X140Y115_DO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D1 = CLBLM_L_X98Y111_SLICE_X155Y111_AQ;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B3 = CLBLL_L_X102Y122_SLICE_X160Y122_C5Q;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D5 = CLBLL_L_X100Y111_SLICE_X156Y111_B5Q;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B4 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D6 = CLBLM_R_X101Y111_SLICE_X158Y111_A5Q;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C5 = CLBLM_L_X90Y114_SLICE_X142Y114_AQ;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C6 = CLBLM_L_X90Y117_SLICE_X143Y117_DO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B5 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C3 = CLBLM_L_X90Y114_SLICE_X142Y114_DO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_C4 = CLBLM_L_X90Y115_SLICE_X142Y115_A5Q;
  assign LIOB33_SING_X0Y99_IOB_X0Y99_T = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D1 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D2 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D3 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D4 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D5 = 1'b1;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_D6 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y115_SLICE_X142Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C6 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A1 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A3 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A4 = CLBLL_L_X100Y115_SLICE_X156Y115_AQ;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A5 = CLBLL_L_X100Y111_SLICE_X157Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_A6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B1 = CLBLM_L_X98Y111_SLICE_X154Y111_B5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B3 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B4 = CLBLL_L_X100Y111_SLICE_X157Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B5 = CLBLL_L_X100Y111_SLICE_X157Y111_C5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_B6 = 1'b1;
  assign LIOB33_X0Y233_IOB_X0Y233_O = 1'b0;
  assign LIOB33_X0Y233_IOB_X0Y234_O = 1'b0;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C1 = CLBLM_R_X101Y111_SLICE_X158Y111_CO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C3 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C4 = CLBLL_L_X100Y113_SLICE_X157Y113_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C5 = CLBLM_L_X98Y111_SLICE_X154Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_C6 = 1'b1;
  assign LIOB33_X0Y233_IOB_X0Y233_T = 1'b1;
  assign LIOB33_X0Y233_IOB_X0Y234_T = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D2 = CLBLM_R_X97Y111_SLICE_X152Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D3 = CLBLM_R_X101Y111_SLICE_X158Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D4 = CLBLM_R_X101Y111_SLICE_X159Y111_B5Q;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_D6 = CLBLL_L_X100Y111_SLICE_X157Y111_AQ;
  assign CLBLL_L_X100Y111_SLICE_X157Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A5 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A6 = 1'b1;
  assign LIOB33_X0Y239_IOB_X0Y240_O = 1'b0;
  assign LIOB33_X0Y239_IOB_X0Y239_O = 1'b0;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A1 = CLBLM_R_X93Y128_SLICE_X147Y128_A5Q;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A2 = CLBLM_R_X93Y128_SLICE_X147Y128_B5Q;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A3 = CLBLM_R_X93Y131_SLICE_X146Y131_A5Q;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A5 = CLBLM_L_X92Y129_SLICE_X145Y129_A5Q;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_A6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B6 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B1 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B2 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B4 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B5 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_B6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_T = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = 1'b0;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C1 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C2 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C4 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C5 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_C6 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C1 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D1 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D2 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D4 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D5 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_D6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C2 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X147Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y239_IOB_X0Y239_T = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C2 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A1 = CLBLM_R_X93Y129_SLICE_X146Y129_BQ;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A4 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C3 = CLBLM_R_X93Y117_SLICE_X146Y117_BQ;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A5 = CLBLM_R_X93Y129_SLICE_X146Y129_A5Q;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_A6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C5 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D4 = CLBLM_R_X89Y119_SLICE_X141Y119_A5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B1 = CLBLM_R_X93Y129_SLICE_X146Y129_B5Q;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B4 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B5 = CLBLM_L_X94Y125_SLICE_X148Y125_A5Q;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_B6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D5 = CLBLM_R_X89Y119_SLICE_X141Y119_AQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D6 = CLBLM_R_X89Y118_SLICE_X141Y118_CQ;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C5 = CLBLM_R_X93Y117_SLICE_X146Y117_B5Q;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_C6 = CLBLM_L_X90Y115_SLICE_X143Y115_BQ;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C2 = CLBLM_R_X95Y130_SLICE_X151Y130_DO6;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C3 = CLBLM_R_X93Y129_SLICE_X146Y129_BQ;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_C6 = CLBLM_R_X93Y126_SLICE_X146Y126_BO6;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D1 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D2 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D3 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D4 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D5 = 1'b1;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_D6 = 1'b1;
  assign CLBLM_R_X93Y117_SLICE_X146Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y129_SLICE_X146Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A1 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A2 = CLBLM_R_X89Y116_SLICE_X140Y116_AQ;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A4 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A5 = CLBLM_L_X90Y116_SLICE_X143Y116_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_A6 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B1 = CLBLM_L_X90Y116_SLICE_X143Y116_DO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B2 = CLBLM_L_X90Y115_SLICE_X143Y115_C5Q;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A4 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B5 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B6 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_B4 = CLBLM_L_X90Y117_SLICE_X143Y117_B5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C2 = CLBLM_L_X90Y116_SLICE_X142Y116_A5Q;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A6 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C3 = CLBLM_L_X92Y116_SLICE_X144Y116_B5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C4 = CLBLM_L_X92Y116_SLICE_X144Y116_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C5 = CLBLM_L_X90Y116_SLICE_X143Y116_CQ;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_C6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A1 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A3 = CLBLL_L_X100Y112_SLICE_X156Y112_AQ;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A4 = CLBLM_L_X98Y112_SLICE_X154Y112_BQ;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A5 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_A6 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D1 = CLBLM_L_X92Y120_SLICE_X144Y120_DO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D2 = CLBLM_L_X90Y116_SLICE_X142Y116_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D4 = CLBLM_R_X89Y114_SLICE_X141Y114_CO6;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_D6 = CLBLM_R_X89Y116_SLICE_X140Y116_AQ;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y116_SLICE_X143Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C2 = CLBLL_L_X100Y112_SLICE_X156Y112_AQ;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B4 = CLBLM_R_X97Y112_SLICE_X152Y112_DO6;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A1 = CLBLM_R_X89Y114_SLICE_X141Y114_B5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A2 = CLBLM_L_X90Y115_SLICE_X142Y115_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A3 = CLBLM_L_X92Y116_SLICE_X145Y116_CO6;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A4 = CLBLM_L_X90Y119_SLICE_X142Y119_C5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_A6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C4 = CLBLL_L_X100Y112_SLICE_X156Y112_A5Q;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C5 = CLBLL_L_X100Y113_SLICE_X156Y113_A5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B1 = CLBLM_L_X90Y117_SLICE_X142Y117_CQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B2 = CLBLM_L_X90Y116_SLICE_X142Y116_BQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B4 = CLBLM_L_X90Y115_SLICE_X142Y115_BQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B5 = CLBLM_L_X90Y116_SLICE_X142Y116_C5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_B6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D1 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D2 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D4 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D5 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_D6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C2 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C3 = CLBLM_L_X90Y116_SLICE_X142Y116_AQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C4 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C5 = CLBLM_L_X90Y117_SLICE_X142Y117_CQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_C6 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B6 = 1'b1;
  assign LIOB33_X0Y235_IOB_X0Y235_O = 1'b0;
  assign LIOB33_X0Y235_IOB_X0Y236_O = 1'b0;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D1 = CLBLM_L_X90Y116_SLICE_X142Y116_C5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D2 = CLBLM_R_X95Y117_SLICE_X150Y117_C5Q;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D4 = CLBLM_L_X90Y116_SLICE_X142Y116_BQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D5 = CLBLM_L_X90Y117_SLICE_X142Y117_CQ;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_D6 = CLBLM_L_X90Y115_SLICE_X142Y115_BQ;
  assign LIOB33_X0Y235_IOB_X0Y235_T = 1'b1;
  assign LIOB33_X0Y235_IOB_X0Y236_T = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A1 = CLBLL_L_X102Y112_SLICE_X160Y112_CO6;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A4 = CLBLM_R_X101Y112_SLICE_X158Y112_B5Q;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A5 = CLBLL_L_X100Y113_SLICE_X156Y113_A5Q;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_A6 = 1'b1;
  assign CLBLM_L_X90Y116_SLICE_X142Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B1 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B2 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B4 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B5 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_B6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C1 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C2 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C1 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C2 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C4 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C5 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_C6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C4 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D1 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D2 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D3 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D4 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D5 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_D6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X157Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = 1'b0;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = 1'b0;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = 1'b0;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_D1 = 1'b0;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_T = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_T1 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A1 = CLBLM_R_X93Y130_SLICE_X147Y130_BO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A2 = CLBLM_R_X95Y130_SLICE_X150Y130_DO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A3 = CLBLM_R_X93Y130_SLICE_X146Y130_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_D1 = 1'b0;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_AX = CLBLM_R_X93Y130_SLICE_X147Y130_BO5;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B1 = CLBLM_R_X93Y130_SLICE_X147Y130_CQ;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B3 = CLBLM_R_X93Y130_SLICE_X147Y130_AQ;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B4 = CLBLM_R_X93Y130_SLICE_X147Y130_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B5 = CLBLM_R_X93Y130_SLICE_X147Y130_C5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = 1'b0;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign RIOB33_X105Y83_IOB_X1Y84_O = CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C2 = CLBLM_R_X93Y130_SLICE_X147Y130_CQ;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C3 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C4 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C5 = CLBLM_R_X93Y130_SLICE_X147Y130_AQ;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_C6 = 1'b1;
  assign RIOB33_X105Y83_IOB_X1Y83_O = CLBLL_L_X102Y117_SLICE_X160Y117_CO6;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D1 = CLBLM_R_X93Y130_SLICE_X147Y130_C5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D2 = CLBLM_R_X93Y130_SLICE_X147Y130_CQ;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D4 = CLBLM_R_X93Y130_SLICE_X147Y130_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D5 = CLBLM_R_X93Y130_SLICE_X147Y130_AQ;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_D6 = CLBLM_L_X92Y131_SLICE_X144Y131_C5Q;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = 1'b0;
  assign CLBLM_R_X93Y130_SLICE_X147Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A1 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A2 = CLBLM_R_X93Y130_SLICE_X146Y130_A5Q;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A3 = CLBLM_R_X93Y132_SLICE_X146Y132_AQ;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A5 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B1 = CLBLM_R_X93Y130_SLICE_X146Y130_B5Q;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B3 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B4 = CLBLM_R_X93Y129_SLICE_X146Y129_AQ;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B5 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C1 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C2 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C3 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C4 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C5 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_C6 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D1 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A2 = CLBLL_L_X100Y112_SLICE_X156Y112_BO6;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D3 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D4 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D5 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_D6 = 1'b1;
  assign CLBLM_R_X93Y130_SLICE_X146Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A1 = CLBLM_R_X93Y119_SLICE_X146Y119_AQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A2 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A4 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A5 = CLBLM_L_X90Y118_SLICE_X143Y118_B5Q;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_A6 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b0;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B1 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B2 = CLBLM_L_X90Y117_SLICE_X143Y117_BQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B4 = CLBLM_L_X90Y117_SLICE_X143Y117_AQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B5 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_B6 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_T = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C1 = CLBLM_L_X90Y116_SLICE_X143Y116_A5Q;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C3 = CLBLM_L_X92Y119_SLICE_X145Y119_DO6;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C4 = CLBLM_L_X90Y116_SLICE_X143Y116_CQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_C6 = CLBLM_L_X90Y118_SLICE_X142Y118_DO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A3 = CLBLL_L_X100Y112_SLICE_X156Y112_A5Q;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A5 = CLBLM_L_X98Y113_SLICE_X154Y113_AQ;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D1 = CLBLM_L_X90Y117_SLICE_X143Y117_BQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D2 = CLBLM_L_X90Y117_SLICE_X143Y117_AQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D4 = CLBLM_R_X93Y119_SLICE_X146Y119_AQ;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D5 = CLBLM_L_X90Y117_SLICE_X143Y117_B5Q;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_D6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B5 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X143Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C1 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C2 = CLBLM_R_X101Y113_SLICE_X158Y113_CO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B6 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A2 = CLBLM_R_X89Y117_SLICE_X140Y117_A5Q;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A3 = CLBLM_R_X89Y116_SLICE_X141Y116_DO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A4 = CLBLM_L_X90Y117_SLICE_X142Y117_BO6;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D1 = CLBLM_L_X98Y113_SLICE_X154Y113_AQ;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D2 = CLBLL_L_X100Y113_SLICE_X156Y113_AQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_AX = CLBLM_L_X90Y117_SLICE_X142Y117_BO5;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D3 = CLBLL_L_X100Y113_SLICE_X156Y113_BQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B1 = CLBLM_L_X90Y117_SLICE_X142Y117_AQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B2 = CLBLM_L_X90Y117_SLICE_X142Y117_A5Q;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D5 = CLBLL_L_X100Y113_SLICE_X156Y113_B5Q;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B4 = CLBLM_L_X90Y119_SLICE_X142Y119_BQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B5 = CLBLM_L_X90Y117_SLICE_X142Y117_C5Q;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_B6 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C1 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C3 = CLBLM_L_X90Y119_SLICE_X142Y119_BQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C4 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C5 = CLBLM_L_X90Y115_SLICE_X142Y115_BQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_C6 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C3 = 1'b1;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D1 = CLBLM_L_X90Y117_SLICE_X142Y117_C5Q;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D2 = CLBLM_L_X90Y117_SLICE_X142Y117_AQ;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D3 = CLBLM_R_X95Y117_SLICE_X150Y117_CQ;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_D6 = CLBLM_L_X90Y119_SLICE_X142Y119_BQ;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A3 = CLBLM_L_X98Y114_SLICE_X154Y114_C5Q;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A4 = CLBLL_L_X100Y113_SLICE_X157Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A5 = CLBLL_L_X100Y115_SLICE_X156Y115_B5Q;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B3 = CLBLM_R_X101Y112_SLICE_X159Y112_DO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B4 = CLBLM_L_X98Y110_SLICE_X154Y110_BO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B5 = CLBLL_L_X100Y115_SLICE_X156Y115_AQ;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B6 = CLBLL_L_X102Y113_SLICE_X161Y113_A5Q;
  assign CLBLM_L_X90Y117_SLICE_X142Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = 1'b0;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C1 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D1 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_SING_X0Y200_IOB_X0Y200_O = 1'b0;
  assign LIOB33_SING_X0Y200_IOB_X0Y200_T = 1'b1;
  assign RIOB33_X105Y85_IOB_X1Y86_O = CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  assign RIOB33_X105Y85_IOB_X1Y85_O = CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A1 = CLBLM_R_X93Y133_SLICE_X146Y133_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A2 = CLBLM_L_X92Y131_SLICE_X145Y131_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A3 = CLBLM_R_X93Y131_SLICE_X147Y131_AQ;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A4 = CLBLM_R_X93Y129_SLICE_X147Y129_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_A6 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B1 = CLBLM_R_X93Y130_SLICE_X147Y130_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B2 = CLBLM_R_X93Y131_SLICE_X147Y131_BQ;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B4 = CLBLM_L_X92Y132_SLICE_X145Y132_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B5 = CLBLM_R_X93Y131_SLICE_X147Y131_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_B6 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C1 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C2 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C3 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C4 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C5 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_C6 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D1 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D2 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D3 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D4 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D5 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_D6 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X147Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A1 = CLBLM_R_X97Y131_SLICE_X152Y131_DO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A4 = CLBLM_R_X93Y131_SLICE_X146Y131_BO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_A6 = CLBLM_R_X93Y130_SLICE_X146Y130_B5Q;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_AX = CLBLM_R_X93Y131_SLICE_X146Y131_BO5;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B1 = CLBLM_R_X93Y131_SLICE_X146Y131_CQ;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B2 = CLBLM_R_X93Y131_SLICE_X146Y131_AQ;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B4 = CLBLM_R_X93Y131_SLICE_X146Y131_A5Q;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B5 = CLBLM_R_X93Y131_SLICE_X146Y131_C5Q;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_B6 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A3 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C2 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C3 = CLBLM_R_X93Y131_SLICE_X146Y131_AQ;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C4 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C5 = CLBLM_R_X93Y131_SLICE_X146Y131_CQ;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_C6 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B5 = CLBLM_L_X98Y112_SLICE_X154Y112_CO6;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D1 = CLBLM_R_X93Y131_SLICE_X146Y131_C5Q;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D2 = CLBLM_R_X93Y131_SLICE_X146Y131_AQ;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D4 = CLBLM_R_X93Y131_SLICE_X146Y131_A5Q;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B6 = 1'b1;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D5 = CLBLM_R_X93Y131_SLICE_X146Y131_CQ;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_D6 = CLBLM_L_X90Y128_SLICE_X143Y128_D5Q;
  assign LIOB33_SING_X0Y249_IOB_X0Y249_T = 1'b1;
  assign LIOB33_SING_X0Y249_IOB_X0Y249_O = 1'b0;
  assign CLBLM_R_X93Y131_SLICE_X146Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A1 = CLBLM_L_X92Y114_SLICE_X145Y114_AQ;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A2 = CLBLM_L_X90Y118_SLICE_X143Y118_A5Q;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A4 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A5 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_A6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B1 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B2 = CLBLM_L_X90Y118_SLICE_X143Y118_BQ;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B4 = CLBLM_R_X93Y119_SLICE_X146Y119_BQ;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A2 = CLBLL_L_X100Y114_SLICE_X156Y114_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A3 = CLBLM_L_X98Y112_SLICE_X154Y112_AQ;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A4 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A5 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_A6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_B6 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B2 = CLBLM_R_X101Y114_SLICE_X158Y114_CO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C4 = CLBLM_L_X98Y112_SLICE_X154Y112_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B3 = CLBLL_L_X100Y113_SLICE_X156Y113_C5Q;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B4 = CLBLM_L_X98Y115_SLICE_X155Y115_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_B6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C6 = CLBLM_R_X97Y113_SLICE_X152Y113_BO6;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D2 = CLBLM_L_X90Y117_SLICE_X143Y117_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C1 = CLBLL_L_X100Y114_SLICE_X156Y114_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C2 = CLBLM_L_X94Y115_SLICE_X148Y115_DO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C4 = CLBLM_L_X98Y115_SLICE_X155Y115_DO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C5 = CLBLL_L_X100Y114_SLICE_X156Y114_B5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D3 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D5 = CLBLM_L_X90Y118_SLICE_X143Y118_B5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D1 = CLBLM_R_X101Y113_SLICE_X159Y113_DO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D2 = CLBLM_L_X98Y114_SLICE_X154Y114_DO6;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D4 = CLBLL_L_X100Y115_SLICE_X156Y115_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D5 = CLBLL_L_X102Y114_SLICE_X160Y114_B5Q;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A5 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A6 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X156Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B1 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B2 = CLBLM_L_X90Y118_SLICE_X142Y118_BQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B4 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B5 = CLBLM_L_X90Y120_SLICE_X143Y120_AQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_B6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C1 = CLBLM_R_X95Y118_SLICE_X150Y118_CQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C2 = CLBLM_R_X89Y118_SLICE_X140Y118_BQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C3 = CLBLM_R_X89Y118_SLICE_X140Y118_B5Q;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C4 = CLBLM_L_X90Y118_SLICE_X142Y118_A5Q;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_C6 = CLBLM_R_X89Y118_SLICE_X140Y118_DQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A1 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A2 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A3 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A4 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A5 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_A6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D1 = CLBLM_L_X90Y120_SLICE_X143Y120_AQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D2 = CLBLM_L_X92Y116_SLICE_X144Y116_A5Q;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B1 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B2 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B3 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B4 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B5 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_B6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C1 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C2 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C3 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C4 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C5 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_C6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C1 = CLBLM_L_X90Y115_SLICE_X143Y115_AQ;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D1 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D2 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D3 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D4 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D5 = 1'b1;
  assign CLBLL_L_X100Y114_SLICE_X157Y114_D6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C4 = CLBLM_L_X92Y116_SLICE_X145Y116_A5Q;
  assign LIOB33_X0Y1_IOB_X0Y1_O = 1'b0;
  assign LIOB33_X0Y1_IOB_X0Y2_O = 1'b0;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C6 = CLBLM_L_X90Y118_SLICE_X142Y118_DO6;
  assign LIOB33_X0Y1_IOB_X0Y2_T = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_T = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A1 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A2 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A3 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A4 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A5 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_A6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B1 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B2 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B3 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B4 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B5 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_B6 = 1'b1;
  assign RIOB33_X105Y87_IOB_X1Y87_O = CLBLL_L_X100Y115_SLICE_X157Y115_CO6;
  assign RIOB33_X105Y87_IOB_X1Y88_O = CLBLM_R_X101Y117_SLICE_X159Y117_AO5;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C1 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C2 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C3 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C4 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C5 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_C6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D1 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D2 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D3 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D4 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D5 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X159Y110_D6 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y4_O = 1'b0;
  assign LIOB33_X0Y3_IOB_X0Y3_O = 1'b0;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A1 = CLBLM_R_X101Y110_SLICE_X158Y110_B5Q;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A2 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A3 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A5 = CLBLL_L_X100Y111_SLICE_X157Y111_BQ;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_A6 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A2 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A3 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D6 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A4 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_A6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B1 = CLBLL_L_X100Y111_SLICE_X157Y111_CQ;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B2 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B4 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_B6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B5 = CLBLM_R_X101Y110_SLICE_X158Y110_BQ;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_B6 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C2 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C4 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_C6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C5 = CLBLM_R_X101Y110_SLICE_X158Y110_B5Q;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_C6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D1 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D2 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D2 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D4 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X147Y132_D6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D4 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D5 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_D6 = 1'b1;
  assign CLBLM_R_X101Y110_SLICE_X158Y110_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A2 = CLBLM_R_X93Y132_SLICE_X146Y132_A5Q;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A3 = CLBLM_R_X93Y130_SLICE_X146Y130_BQ;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = 1'b0;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B2 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B4 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B5 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A6 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C2 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C4 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = 1'b0;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C1 = CLBLM_L_X90Y115_SLICE_X143Y115_C5Q;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D1 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D2 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C3 = CLBLM_R_X93Y119_SLICE_X146Y119_DO6;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D3 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D4 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D5 = 1'b1;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_D6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C4 = CLBLM_L_X90Y118_SLICE_X143Y118_A5Q;
  assign LIOB33_X0Y241_IOB_X0Y242_O = 1'b0;
  assign CLBLM_R_X93Y132_SLICE_X146Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y241_IOB_X0Y241_O = 1'b0;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_D1 = 1'b0;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_C6 = CLBLM_L_X90Y118_SLICE_X143Y118_DO6;
  assign LIOB33_X0Y241_IOB_X0Y242_T = 1'b1;
  assign LIOB33_X0Y241_IOB_X0Y241_T = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_T1 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A1 = CLBLM_L_X90Y119_SLICE_X143Y119_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A2 = CLBLM_L_X90Y120_SLICE_X143Y120_BQ;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A4 = CLBLM_L_X90Y119_SLICE_X143Y119_CQ;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A5 = CLBLM_L_X90Y120_SLICE_X143Y120_CQ;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_A6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A2 = CLBLL_L_X100Y115_SLICE_X156Y115_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A3 = CLBLL_L_X100Y116_SLICE_X156Y116_AQ;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A4 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A5 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_A6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B3 = CLBLL_L_X102Y124_SLICE_X161Y124_DO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_AX = CLBLM_L_X90Y119_SLICE_X142Y119_AO5;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B1 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B2 = CLBLL_L_X100Y114_SLICE_X156Y114_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B3 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B4 = CLBLM_L_X98Y114_SLICE_X154Y114_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C4 = CLBLM_L_X90Y119_SLICE_X142Y119_C5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B5 = CLBLL_L_X100Y115_SLICE_X156Y115_C5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_B6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C1 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C2 = CLBLM_L_X98Y116_SLICE_X155Y116_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C4 = CLBLM_R_X97Y115_SLICE_X153Y115_B5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C5 = CLBLL_L_X100Y115_SLICE_X156Y115_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_C6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_CX = CLBLM_L_X90Y119_SLICE_X143Y119_AO5;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D3 = CLBLM_L_X90Y118_SLICE_X143Y118_AQ;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D4 = CLBLM_L_X94Y124_SLICE_X148Y124_DO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D5 = CLBLM_L_X90Y117_SLICE_X143Y117_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D2 = CLBLM_L_X90Y116_SLICE_X143Y116_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D1 = CLBLL_L_X100Y116_SLICE_X156Y116_AQ;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D2 = CLBLL_L_X102Y115_SLICE_X160Y115_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D3 = CLBLM_L_X98Y115_SLICE_X154Y115_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D5 = CLBLM_R_X101Y116_SLICE_X158Y116_DO6;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y115_SLICE_X156Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C1 = CLBLL_L_X102Y123_SLICE_X160Y123_AQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A1 = CLBLM_L_X90Y119_SLICE_X142Y119_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A2 = CLBLM_R_X89Y117_SLICE_X140Y117_BQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C2 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D4 = CLBLM_L_X90Y118_SLICE_X143Y118_BQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A5 = CLBLM_L_X90Y119_SLICE_X143Y119_AQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B1 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C3 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B2 = CLBLM_L_X90Y118_SLICE_X142Y118_AQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y118_SLICE_X143Y118_D6 = CLBLM_R_X93Y119_SLICE_X146Y119_BQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C2 = CLBLM_R_X89Y120_SLICE_X141Y120_C5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C3 = CLBLM_R_X89Y115_SLICE_X140Y115_A5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C4 = CLBLM_R_X89Y116_SLICE_X140Y116_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C5 = CLBLM_L_X90Y119_SLICE_X142Y119_CQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_C6 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A3 = CLBLM_L_X98Y117_SLICE_X154Y117_AO6;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A4 = CLBLL_L_X100Y115_SLICE_X157Y115_DO6;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_A6 = CLBLL_L_X102Y117_SLICE_X161Y117_A5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D3 = CLBLM_L_X90Y118_SLICE_X142Y118_AQ;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D5 = CLBLM_L_X90Y119_SLICE_X142Y119_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D6 = CLBLM_R_X89Y117_SLICE_X140Y117_BQ;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B2 = CLBLL_L_X100Y115_SLICE_X157Y115_BQ;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B3 = CLBLL_L_X100Y115_SLICE_X157Y115_AQ;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B4 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B5 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_B6 = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C1 = CLBLL_L_X100Y115_SLICE_X157Y115_BQ;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C2 = CLBLL_L_X100Y115_SLICE_X157Y115_AQ;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C3 = CLBLM_R_X101Y115_SLICE_X158Y115_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C4 = CLBLL_L_X102Y117_SLICE_X161Y117_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C5 = CLBLL_L_X100Y115_SLICE_X157Y115_B5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A2 = CLBLM_L_X98Y133_SLICE_X154Y133_BQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A1 = CLBLM_R_X89Y118_SLICE_X140Y118_DQ;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A3 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y3_T = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y4_T = 1'b1;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D1 = CLBLL_L_X100Y115_SLICE_X157Y115_BQ;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D2 = CLBLM_R_X101Y115_SLICE_X158Y115_A5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D4 = CLBLL_L_X100Y115_SLICE_X157Y115_AQ;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D5 = CLBLL_L_X100Y115_SLICE_X157Y115_B5Q;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_D6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A2 = CLBLM_R_X89Y117_SLICE_X140Y117_BQ;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y115_SLICE_X157Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_A4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A5 = CLBLM_L_X98Y133_SLICE_X154Y133_A5Q;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D1 = CLBLL_L_X102Y124_SLICE_X160Y124_DQ;
  assign RIOB33_X105Y89_IOB_X1Y90_O = CLBLL_L_X102Y116_SLICE_X160Y116_AO6;
  assign RIOB33_X105Y89_IOB_X1Y89_O = CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D2 = CLBLL_L_X102Y124_SLICE_X161Y124_A5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D3 = CLBLM_L_X92Y116_SLICE_X144Y116_BQ;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D3 = CLBLL_L_X102Y124_SLICE_X161Y124_B5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D4 = CLBLM_L_X92Y119_SLICE_X144Y119_CQ;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D5 = CLBLM_L_X92Y116_SLICE_X144Y116_B5Q;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D5 = CLBLL_L_X102Y120_SLICE_X160Y120_D5Q;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A1 = CLBLM_R_X101Y111_SLICE_X159Y111_B5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A2 = CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A3 = CLBLM_R_X101Y111_SLICE_X158Y111_A5Q;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_D6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A5 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_A6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B2 = CLBLM_L_X98Y133_SLICE_X154Y133_B5Q;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B1 = CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B2 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B3 = CLBLL_L_X102Y111_SLICE_X161Y111_DO6;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B3 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B5 = CLBLM_R_X101Y111_SLICE_X158Y111_B5Q;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_B6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B4 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C1 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C2 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C3 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B5 = CLBLM_L_X98Y133_SLICE_X155Y133_AQ;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C4 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C5 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_C6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_B6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D1 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D2 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D3 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D4 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D5 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_D6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X159Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A1 = CLBLM_L_X98Y112_SLICE_X155Y112_AQ;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A2 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A3 = CLBLL_L_X100Y111_SLICE_X156Y111_B5Q;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A5 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_A6 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A1 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A3 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C1 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A5 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_A6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B1 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B3 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C3 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B5 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_B6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_B6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C4 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C1 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C3 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C5 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C5 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_C6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C5 = CLBLL_L_X100Y111_SLICE_X157Y111_A5Q;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_C6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D1 = CLBLM_R_X101Y110_SLICE_X158Y110_AQ;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D1 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D3 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D4 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D5 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X147Y133_D6 = 1'b1;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D3 = CLBLM_R_X101Y111_SLICE_X158Y111_BQ;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D4 = CLBLL_L_X100Y111_SLICE_X157Y111_BQ;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y111_SLICE_X158Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A3 = CLBLM_R_X93Y132_SLICE_X146Y132_A5Q;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A4 = CLBLM_R_X93Y133_SLICE_X146Y133_BO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_A6 = CLBLM_L_X94Y132_SLICE_X149Y132_AO6;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_AX = CLBLM_R_X93Y133_SLICE_X146Y133_BO5;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B1 = CLBLM_R_X93Y133_SLICE_X146Y133_CQ;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B2 = CLBLM_R_X93Y133_SLICE_X146Y133_C5Q;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B3 = CLBLM_R_X93Y133_SLICE_X146Y133_AQ;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B4 = CLBLM_R_X93Y133_SLICE_X146Y133_A5Q;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_B6 = 1'b1;
  assign LIOB33_X0Y243_IOB_X0Y243_O = 1'b0;
  assign LIOB33_X0Y243_IOB_X0Y244_O = 1'b0;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C3 = CLBLM_R_X93Y133_SLICE_X146Y133_AQ;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C4 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C5 = CLBLM_R_X93Y133_SLICE_X146Y133_CQ;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_C6 = 1'b1;
  assign LIOB33_X0Y243_IOB_X0Y243_T = 1'b1;
  assign LIOB33_X0Y243_IOB_X0Y244_T = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D1 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D1 = CLBLM_R_X93Y133_SLICE_X146Y133_C5Q;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D3 = CLBLM_R_X93Y133_SLICE_X146Y133_AQ;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D2 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D4 = CLBLM_R_X93Y133_SLICE_X146Y133_A5Q;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D5 = CLBLM_R_X93Y133_SLICE_X146Y133_CQ;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_D6 = CLBLM_L_X92Y131_SLICE_X144Y131_B5Q;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D3 = 1'b1;
  assign CLBLM_R_X93Y133_SLICE_X146Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D4 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D3 = CLBLM_L_X90Y118_SLICE_X142Y118_BQ;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D6 = 1'b1;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D4 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A2 = CLBLM_L_X90Y117_SLICE_X143Y117_CO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A2 = CLBLL_L_X100Y116_SLICE_X156Y116_A5Q;
  assign CLBLM_L_X90Y118_SLICE_X142Y118_D5 = CLBLM_L_X90Y118_SLICE_X142Y118_B5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A3 = CLBLL_L_X100Y117_SLICE_X157Y117_AQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A4 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A5 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_A6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A3 = CLBLM_L_X92Y122_SLICE_X144Y122_C5Q;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A5 = CLBLM_L_X90Y122_SLICE_X143Y122_C5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B2 = CLBLL_L_X100Y116_SLICE_X156Y116_BQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B3 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B4 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B5 = CLBLM_L_X98Y116_SLICE_X155Y116_AQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_B6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B5 = CLBLM_L_X90Y120_SLICE_X142Y120_AQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C1 = CLBLM_R_X97Y115_SLICE_X153Y115_DO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C3 = CLBLL_L_X102Y116_SLICE_X160Y116_B5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C4 = CLBLL_L_X100Y116_SLICE_X156Y116_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C5 = CLBLL_L_X100Y116_SLICE_X156Y116_DO6;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C2 = CLBLM_R_X89Y120_SLICE_X141Y120_AQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D1 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D2 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D1 = CLBLM_L_X98Y116_SLICE_X155Y116_AQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D2 = CLBLM_R_X101Y116_SLICE_X158Y116_A5Q;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D3 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D4 = CLBLL_L_X100Y116_SLICE_X156Y116_BQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D5 = CLBLL_L_X100Y116_SLICE_X156Y116_B5Q;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B2 = CLBLL_L_X102Y124_SLICE_X161Y124_BQ;
  assign CLBLL_L_X100Y116_SLICE_X156Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A1 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A2 = CLBLM_L_X90Y120_SLICE_X142Y120_A5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A4 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A5 = CLBLM_R_X89Y122_SLICE_X141Y122_AQ;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_A6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B1 = CLBLM_R_X93Y124_SLICE_X146Y124_DO6;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B5 = CLBLM_L_X90Y120_SLICE_X142Y120_A5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_B6 = CLBLM_L_X90Y120_SLICE_X142Y120_CO6;
  assign LIOB33_X0Y5_IOB_X0Y5_O = 1'b0;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B6 = 1'b1;
  assign LIOB33_X0Y5_IOB_X0Y6_O = 1'b0;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_BX = CLBLM_L_X90Y120_SLICE_X142Y120_CO5;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C1 = CLBLM_L_X90Y120_SLICE_X142Y120_BQ;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C2 = CLBLM_R_X89Y120_SLICE_X141Y120_AQ;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C3 = CLBLM_L_X90Y120_SLICE_X143Y120_C5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A2 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A3 = CLBLL_L_X100Y116_SLICE_X157Y116_AQ;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A4 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A5 = CLBLM_L_X98Y115_SLICE_X155Y115_AQ;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_A6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C5 = CLBLM_L_X90Y120_SLICE_X142Y120_B5Q;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_C6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B2 = CLBLL_L_X100Y116_SLICE_X157Y116_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B3 = CLBLL_L_X100Y114_SLICE_X156Y114_B5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B4 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D3 = CLBLM_L_X90Y120_SLICE_X143Y120_C5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B5 = CLBLM_R_X101Y116_SLICE_X158Y116_CO6;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D4 = CLBLM_L_X90Y119_SLICE_X142Y119_CQ;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D5 = CLBLM_L_X90Y120_SLICE_X142Y120_B5Q;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_B6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D1 = CLBLM_L_X90Y120_SLICE_X142Y120_BQ;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C2 = CLBLL_L_X102Y124_SLICE_X160Y124_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C2 = CLBLL_L_X100Y117_SLICE_X157Y117_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C4 = CLBLL_L_X100Y118_SLICE_X156Y118_CO6;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C3 = CLBLL_L_X102Y124_SLICE_X161Y124_BQ;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C5 = CLBLL_L_X100Y117_SLICE_X157Y117_B5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_C6 = CLBLM_L_X92Y116_SLICE_X145Y116_DO6;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C4 = CLBLM_R_X95Y116_SLICE_X150Y116_A5Q;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C5 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D1 = CLBLM_L_X98Y115_SLICE_X155Y115_AQ;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D2 = 1'b1;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D4 = CLBLL_L_X100Y116_SLICE_X157Y116_A5Q;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D5 = CLBLL_L_X100Y116_SLICE_X157Y116_AQ;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_D6 = CLBLM_R_X97Y115_SLICE_X152Y115_AQ;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C6 = CLBLM_R_X95Y115_SLICE_X150Y115_A5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y116_SLICE_X157Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_T1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A1 = CLBLL_L_X100Y113_SLICE_X157Y113_AQ;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A2 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A3 = CLBLM_R_X101Y113_SLICE_X159Y113_C5Q;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A5 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_A6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A5 = CLBLM_R_X101Y133_SLICE_X159Y133_AQ;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B3 = CLBLM_R_X101Y112_SLICE_X159Y112_AQ;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B4 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B5 = CLBLM_R_X101Y112_SLICE_X159Y112_BQ;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_B6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A6 = CLBLM_R_X101Y133_SLICE_X158Y133_CO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D2 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C2 = CLBLL_L_X100Y112_SLICE_X157Y112_AQ;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C3 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D3 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C5 = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_C6 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D4 = CLBLL_L_X102Y124_SLICE_X161Y124_AQ;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D5 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D1 = CLBLM_R_X101Y112_SLICE_X159Y112_BQ;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D2 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D4 = CLBLL_L_X100Y113_SLICE_X157Y113_AQ;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D5 = CLBLM_R_X101Y112_SLICE_X159Y112_B5Q;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_D6 = CLBLM_R_X101Y112_SLICE_X159Y112_AQ;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_D1 = 1'b0;
  assign CLBLM_R_X101Y112_SLICE_X159Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A2 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A3 = CLBLM_R_X101Y112_SLICE_X158Y112_AQ;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A5 = CLBLM_R_X101Y111_SLICE_X158Y111_AQ;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_A6 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B2 = CLBLM_R_X101Y112_SLICE_X158Y112_A5Q;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B3 = CLBLM_R_X101Y111_SLICE_X159Y111_A5Q;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B5 = CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_B6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B6 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C1 = CLBLM_R_X101Y111_SLICE_X158Y111_AQ;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C2 = CLBLM_R_X101Y112_SLICE_X158Y112_AQ;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C3 = CLBLM_L_X98Y112_SLICE_X155Y112_AQ;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C4 = CLBLM_R_X101Y112_SLICE_X158Y112_A5Q;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_C6 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D1 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D2 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D3 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D4 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B6 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D5 = 1'b1;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_D6 = 1'b1;
  assign LIOB33_X0Y245_IOB_X0Y245_O = 1'b0;
  assign LIOB33_X0Y245_IOB_X0Y246_O = 1'b0;
  assign CLBLM_R_X101Y112_SLICE_X158Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C1 = CLBLM_R_X101Y130_SLICE_X158Y130_AQ;
  assign LIOB33_X0Y245_IOB_X0Y246_T = 1'b1;
  assign LIOB33_X0Y245_IOB_X0Y245_T = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C2 = CLBLM_R_X101Y133_SLICE_X158Y133_AQ;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y213_T1 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D2 = CLBLM_R_X89Y121_SLICE_X141Y121_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D3 = CLBLM_R_X89Y121_SLICE_X141Y121_CQ;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C5 = CLBLM_R_X101Y133_SLICE_X158Y133_B5Q;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C6 = CLBLM_R_X101Y134_SLICE_X158Y134_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D6 = CLBLM_R_X89Y121_SLICE_X141Y121_AQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_D1 = 1'b0;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A1 = CLBLM_R_X89Y125_SLICE_X141Y125_DO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A3 = CLBLM_L_X90Y121_SLICE_X142Y121_A5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A5 = CLBLL_L_X100Y117_SLICE_X156Y117_CO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A6 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A4 = CLBLM_L_X90Y121_SLICE_X143Y121_BO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A1 = CLBLM_R_X89Y121_SLICE_X140Y121_DO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A2 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_A3 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B3 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B4 = CLBLL_L_X100Y118_SLICE_X156Y118_AQ;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B5 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_B6 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_AX = CLBLM_L_X90Y121_SLICE_X143Y121_BO5;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B1 = CLBLM_L_X90Y121_SLICE_X143Y121_AQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B2 = CLBLM_L_X90Y121_SLICE_X143Y121_A5Q;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B3 = CLBLM_L_X90Y121_SLICE_X143Y121_CQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B5 = CLBLM_L_X90Y121_SLICE_X143Y121_C5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A4 = CLBLM_R_X89Y120_SLICE_X140Y120_BO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C5 = CLBLL_L_X100Y117_SLICE_X156Y117_DO6;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_C6 = CLBLM_L_X98Y116_SLICE_X155Y116_DO6;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C2 = CLBLM_L_X90Y121_SLICE_X143Y121_CQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C3 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C4 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C5 = CLBLM_L_X90Y121_SLICE_X143Y121_AQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_C6 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D2 = CLBLL_L_X100Y117_SLICE_X156Y117_AQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D2 = CLBLM_L_X90Y121_SLICE_X143Y121_CQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D4 = CLBLM_L_X90Y121_SLICE_X143Y121_A5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D3 = CLBLL_L_X100Y117_SLICE_X156Y117_BQ;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D4 = CLBLL_L_X100Y118_SLICE_X156Y118_AQ;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D5 = CLBLL_L_X100Y117_SLICE_X156Y117_B5Q;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_D6 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D1 = CLBLM_L_X90Y121_SLICE_X143Y121_C5Q;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D5 = CLBLM_L_X90Y121_SLICE_X143Y121_AQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_D6 = CLBLM_L_X92Y121_SLICE_X145Y121_CQ;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y117_SLICE_X156Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A1 = CLBLM_L_X90Y114_SLICE_X142Y114_A5Q;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A2 = CLBLM_L_X90Y121_SLICE_X142Y121_A5Q;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A4 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A5 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = 1'b0;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B1 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B2 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B3 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B4 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B5 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_B6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C1 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C2 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C3 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C4 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C5 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_C6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A2 = CLBLM_R_X97Y117_SLICE_X153Y117_AQ;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A3 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A4 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A5 = CLBLL_L_X100Y117_SLICE_X157Y117_A5Q;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_A6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B2 = CLBLM_R_X101Y117_SLICE_X158Y117_CO6;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B3 = CLBLM_R_X97Y117_SLICE_X152Y117_BQ;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B4 = CLBLL_L_X100Y118_SLICE_X156Y118_A5Q;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D2 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D3 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D4 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D5 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B5 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_B6 = 1'b1;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_D1 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C1 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C2 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C3 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C4 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C5 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_C6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y121_SLICE_X142Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D1 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D2 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D3 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D4 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D5 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_D6 = 1'b1;
  assign CLBLL_L_X100Y117_SLICE_X157Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_T1 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C2 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_D1 = 1'b0;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C3 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C4 = CLBLM_R_X89Y120_SLICE_X140Y120_A5Q;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_T1 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C5 = CLBLM_L_X92Y123_SLICE_X144Y123_D5Q;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_C6 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A3 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A4 = CLBLM_R_X101Y113_SLICE_X158Y113_DO6;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A5 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_A6 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_AX = CLBLM_R_X101Y113_SLICE_X159Y113_BO5;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B1 = CLBLM_R_X101Y114_SLICE_X158Y114_DO6;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B3 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B5 = CLBLM_R_X101Y113_SLICE_X159Y113_BQ;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_B6 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_BX = CLBLM_R_X101Y113_SLICE_X159Y113_AO5;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C1 = CLBLL_L_X100Y115_SLICE_X156Y115_BQ;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C2 = CLBLM_R_X101Y113_SLICE_X159Y113_CQ;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C3 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C5 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_C6 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D1 = CLBLL_L_X100Y115_SLICE_X156Y115_BQ;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D2 = CLBLM_R_X101Y113_SLICE_X159Y113_CQ;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D3 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D5 = CLBLM_R_X101Y113_SLICE_X159Y113_C5Q;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_D6 = CLBLM_R_X101Y112_SLICE_X159Y112_A5Q;
  assign CLBLM_R_X101Y113_SLICE_X159Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A1 = CLBLM_R_X101Y113_SLICE_X158Y113_B5Q;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A2 = CLBLL_L_X100Y114_SLICE_X156Y114_BQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A3 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A5 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_A6 = 1'b1;
  assign LIOB33_X0Y247_IOB_X0Y247_O = 1'b0;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B1 = CLBLL_L_X100Y113_SLICE_X156Y113_CQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B3 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B4 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B5 = CLBLM_R_X101Y113_SLICE_X158Y113_BQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_B6 = 1'b1;
  assign LIOB33_X0Y247_IOB_X0Y248_O = 1'b0;
  assign LIOB33_X0Y247_IOB_X0Y248_T = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C1 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C2 = CLBLL_L_X102Y113_SLICE_X160Y113_A5Q;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D6 = CLBLM_R_X97Y120_SLICE_X152Y120_BQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C5 = CLBLM_R_X101Y113_SLICE_X158Y113_DO6;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_C6 = CLBLL_L_X100Y113_SLICE_X156Y113_DO6;
  assign LIOB33_X0Y247_IOB_X0Y247_T = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D1 = CLBLM_R_X101Y113_SLICE_X158Y113_BQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D3 = CLBLL_L_X100Y113_SLICE_X156Y113_CQ;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D4 = CLBLM_R_X101Y113_SLICE_X158Y113_A5Q;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D5 = CLBLM_R_X101Y113_SLICE_X158Y113_B5Q;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_D6 = 1'b1;
  assign CLBLM_R_X101Y113_SLICE_X158Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A2 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A3 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A4 = CLBLL_L_X100Y118_SLICE_X156Y118_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A5 = CLBLL_L_X100Y117_SLICE_X156Y117_AQ;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_A6 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A1 = CLBLM_R_X93Y128_SLICE_X146Y128_DO6;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A4 = CLBLM_L_X90Y122_SLICE_X143Y122_BO6;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A6 = CLBLM_R_X89Y124_SLICE_X141Y124_AQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B2 = CLBLL_L_X100Y118_SLICE_X156Y118_BQ;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B3 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_AX = CLBLM_L_X90Y122_SLICE_X143Y122_BO5;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B2 = CLBLM_L_X90Y124_SLICE_X143Y124_B5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B4 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B5 = CLBLM_L_X90Y122_SLICE_X143Y122_A5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B6 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B1 = CLBLM_L_X90Y122_SLICE_X143Y122_AQ;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_B5 = CLBLM_L_X92Y116_SLICE_X145Y116_AQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_B4 = CLBLM_L_X90Y122_SLICE_X143Y122_CQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C2 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C1 = CLBLL_L_X100Y118_SLICE_X156Y118_BQ;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C2 = CLBLM_L_X92Y116_SLICE_X145Y116_AQ;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C4 = CLBLL_L_X100Y118_SLICE_X156Y118_A5Q;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_C5 = CLBLL_L_X100Y118_SLICE_X156Y118_B5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C3 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C4 = CLBLM_L_X92Y120_SLICE_X144Y120_B5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C5 = CLBLM_L_X90Y122_SLICE_X143Y122_AQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D1 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D2 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D3 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D4 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D5 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_D6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X156Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D1 = CLBLM_R_X89Y120_SLICE_X141Y120_BQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D2 = CLBLM_L_X90Y122_SLICE_X143Y122_CQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D3 = CLBLM_L_X90Y124_SLICE_X143Y124_B5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D4 = CLBLM_L_X90Y122_SLICE_X143Y122_A5Q;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D5 = CLBLM_L_X90Y122_SLICE_X143Y122_AQ;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A1 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A2 = CLBLM_L_X90Y122_SLICE_X142Y122_A5Q;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A4 = CLBLM_L_X90Y121_SLICE_X142Y121_AQ;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A5 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_A6 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B1 = CLBLM_L_X90Y128_SLICE_X142Y128_DO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B2 = CLBLM_L_X92Y122_SLICE_X144Y122_AO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B5 = CLBLM_L_X90Y122_SLICE_X142Y122_A5Q;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_B6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A2 = CLBLM_L_X98Y119_SLICE_X155Y119_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A3 = CLBLL_L_X100Y116_SLICE_X157Y116_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A4 = CLBLM_R_X101Y118_SLICE_X159Y118_CO6;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C1 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C2 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A5 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C4 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C5 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_A6 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_C3 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B2 = CLBLL_L_X100Y118_SLICE_X157Y118_BQ;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B3 = CLBLM_R_X101Y119_SLICE_X159Y119_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B4 = CLBLM_R_X101Y118_SLICE_X158Y118_CQ;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_B5 = CLBLL_L_X102Y117_SLICE_X161Y117_D5Q;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D1 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D2 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D3 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D4 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D5 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_D6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C1 = CLBLM_R_X103Y117_SLICE_X162Y117_B5Q;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C2 = CLBLL_L_X100Y118_SLICE_X157Y118_CQ;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y122_SLICE_X142Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_C6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D1 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D2 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D3 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D4 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D5 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_D6 = 1'b1;
  assign CLBLL_L_X100Y118_SLICE_X157Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A1 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A2 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A3 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A4 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A5 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_A6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B1 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B2 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B3 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B4 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B5 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C1 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C2 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C3 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C4 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C5 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_C6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D1 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D2 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_A6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D3 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D4 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D5 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X159Y114_D6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A1 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A2 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A3 = CLBLM_R_X101Y114_SLICE_X158Y114_AQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A5 = CLBLM_R_X101Y113_SLICE_X158Y113_AQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_A6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B1 = CLBLM_R_X101Y118_SLICE_X159Y118_A5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B2 = CLBLM_R_X101Y114_SLICE_X158Y114_BQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B3 = CLBLL_L_X102Y113_SLICE_X160Y113_A5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B5 = CLBLM_R_X101Y114_SLICE_X158Y114_A5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C1 = CLBLM_R_X101Y114_SLICE_X158Y114_BQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C3 = CLBLM_L_X98Y115_SLICE_X155Y115_DO6;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C5 = CLBLM_R_X101Y114_SLICE_X158Y114_DO6;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_C6 = CLBLM_R_X101Y113_SLICE_X159Y113_BQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D1 = CLBLM_R_X101Y113_SLICE_X158Y113_AQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D2 = 1'b1;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D3 = CLBLM_R_X101Y114_SLICE_X158Y114_AQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D4 = CLBLM_R_X101Y114_SLICE_X158Y114_A5Q;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_D6 = CLBLL_L_X100Y114_SLICE_X156Y114_BQ;
  assign CLBLM_R_X101Y114_SLICE_X158Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D5 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A2 = CLBLL_L_X100Y119_SLICE_X156Y119_B5Q;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A3 = CLBLL_L_X100Y119_SLICE_X156Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A4 = CLBLM_L_X98Y119_SLICE_X155Y119_BQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A5 = CLBLM_L_X98Y119_SLICE_X155Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_A6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B2 = CLBLM_L_X98Y119_SLICE_X155Y119_BQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B3 = CLBLL_L_X100Y120_SLICE_X156Y120_AQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B4 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A4 = CLBLM_L_X90Y123_SLICE_X143Y123_BO6;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A6 = CLBLM_L_X90Y124_SLICE_X143Y124_DO6;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B5 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_B6 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_AX = CLBLM_L_X90Y123_SLICE_X143Y123_BO5;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B1 = CLBLM_L_X90Y123_SLICE_X143Y123_AQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B2 = CLBLM_L_X90Y123_SLICE_X143Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C1 = CLBLM_L_X98Y119_SLICE_X155Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C2 = CLBLL_L_X100Y119_SLICE_X156Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C4 = CLBLM_R_X101Y118_SLICE_X158Y118_CQ;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C5 = CLBLL_L_X100Y119_SLICE_X156Y119_B5Q;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_C6 = CLBLM_L_X98Y119_SLICE_X155Y119_BQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B4 = CLBLM_L_X90Y123_SLICE_X143Y123_CQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C3 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C4 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C5 = CLBLM_L_X90Y123_SLICE_X143Y123_AQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C6 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D1 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D2 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D3 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D4 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D5 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_D6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X156Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D1 = CLBLM_L_X90Y123_SLICE_X143Y123_C5Q;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D2 = CLBLM_L_X90Y123_SLICE_X143Y123_CQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D4 = CLBLM_L_X90Y123_SLICE_X143Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D5 = CLBLM_L_X90Y123_SLICE_X143Y123_AQ;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_D6 = CLBLM_L_X92Y121_SLICE_X144Y121_D5Q;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A1 = CLBLM_L_X90Y122_SLICE_X142Y122_AQ;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A2 = CLBLM_L_X90Y123_SLICE_X142Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A4 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A5 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_A6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A3 = CLBLM_L_X92Y120_SLICE_X145Y120_DO6;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B4 = CLBLM_L_X90Y123_SLICE_X143Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B5 = CLBLM_L_X92Y121_SLICE_X145Y121_AQ;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A4 = CLBLL_L_X100Y119_SLICE_X157Y119_BO6;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_A6 = CLBLM_L_X98Y117_SLICE_X155Y117_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C2 = CLBLM_L_X90Y124_SLICE_X142Y124_A5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_AX = CLBLL_L_X100Y119_SLICE_X157Y119_BO5;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C3 = CLBLM_R_X89Y123_SLICE_X141Y123_A5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C4 = CLBLM_L_X92Y122_SLICE_X144Y122_AQ;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C5 = CLBLM_L_X90Y123_SLICE_X142Y123_B5Q;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_C6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B2 = CLBLM_R_X101Y119_SLICE_X158Y119_A5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B3 = CLBLL_L_X100Y119_SLICE_X157Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B4 = CLBLL_L_X100Y119_SLICE_X157Y119_CQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B5 = CLBLL_L_X100Y119_SLICE_X157Y119_A5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_B6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C1 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C2 = CLBLL_L_X100Y119_SLICE_X156Y119_BQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C4 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C5 = CLBLL_L_X100Y119_SLICE_X157Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_C6 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D6 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D5 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D1 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D2 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D3 = 1'b1;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D1 = CLBLL_L_X100Y119_SLICE_X157Y119_A5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D3 = CLBLL_L_X102Y120_SLICE_X160Y120_BQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D4 = CLBLM_R_X101Y119_SLICE_X158Y119_A5Q;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D5 = CLBLL_L_X100Y119_SLICE_X157Y119_AQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_D6 = CLBLL_L_X100Y119_SLICE_X157Y119_CQ;
  assign CLBLL_L_X100Y119_SLICE_X157Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y5_IOB_X0Y5_T = 1'b1;
  assign LIOB33_X0Y5_IOB_X0Y6_T = 1'b1;
  assign LIOB33_X0Y53_IOB_X0Y54_O = 1'b0;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A2 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A3 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A5 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_A6 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B2 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B3 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B5 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = 1'b0;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C2 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C3 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C5 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_C6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = 1'b0;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D2 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D3 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D5 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X159Y115_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = 1'b0;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A3 = CLBLL_L_X100Y117_SLICE_X157Y117_BQ;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A5 = CLBLL_L_X100Y115_SLICE_X157Y115_B5Q;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = 1'b0;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B3 = CLBLM_R_X101Y115_SLICE_X158Y115_AQ;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B5 = CLBLM_R_X101Y115_SLICE_X158Y115_BQ;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_B6 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_D1 = 1'b0;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C1 = CLBLL_L_X100Y117_SLICE_X157Y117_BQ;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C2 = CLBLM_R_X101Y115_SLICE_X158Y115_AQ;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C3 = CLBLM_R_X101Y115_SLICE_X158Y115_BQ;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C5 = CLBLM_R_X101Y115_SLICE_X158Y115_B5Q;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_C6 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_T1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D1 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D2 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D3 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D4 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D5 = 1'b1;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_D6 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_D1 = 1'b0;
  assign CLBLM_R_X101Y115_SLICE_X158Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B2 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_T1 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B4 = CLBLM_L_X90Y120_SLICE_X143Y120_CQ;
  assign RIOB33_X105Y81_IOB_X1Y82_O = CLBLM_R_X101Y120_SLICE_X159Y120_CO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B5 = CLBLM_R_X93Y124_SLICE_X147Y124_AQ;
  assign RIOB33_X105Y81_IOB_X1Y81_O = CLBLL_L_X102Y119_SLICE_X161Y119_CO6;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_B6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D3 = 1'b1;
  assign RIOB33_X105Y101_IOB_X1Y102_O = 1'b0;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C1 = CLBLM_L_X90Y120_SLICE_X143Y120_CQ;
  assign RIOB33_X105Y101_IOB_X1Y101_O = 1'b0;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C2 = CLBLM_L_X90Y119_SLICE_X143Y119_CQ;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A2 = CLBLL_L_X100Y120_SLICE_X157Y120_BO6;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A5 = CLBLL_L_X100Y121_SLICE_X156Y121_AQ;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_A6 = CLBLM_L_X92Y119_SLICE_X145Y119_CO6;
  assign RIOB33_X105Y101_IOB_X1Y101_T = 1'b1;
  assign RIOB33_X105Y101_IOB_X1Y102_T = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B1 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B2 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B3 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B4 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B5 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_B6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C5 = CLBLM_L_X90Y119_SLICE_X143Y119_B5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A1 = CLBLM_L_X90Y125_SLICE_X142Y125_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A2 = CLBLM_L_X90Y128_SLICE_X143Y128_BQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C1 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C2 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C3 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C4 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A4 = CLBLM_L_X90Y124_SLICE_X143Y124_AQ;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C6 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A5 = CLBLM_L_X90Y124_SLICE_X143Y124_BQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_A6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X143Y119_C6 = CLBLM_L_X90Y120_SLICE_X143Y120_BQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B1 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B2 = CLBLM_L_X90Y122_SLICE_X143Y122_CQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B4 = CLBLM_L_X90Y128_SLICE_X143Y128_BQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B6 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_B5 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D1 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D2 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D3 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D4 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D5 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_D6 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C3 = CLBLM_R_X89Y121_SLICE_X141Y121_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C4 = CLBLM_R_X89Y122_SLICE_X141Y122_B5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C5 = CLBLM_L_X90Y125_SLICE_X143Y125_DQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C6 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D1 = CLBLM_L_X90Y124_SLICE_X143Y124_BQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D2 = CLBLM_L_X90Y124_SLICE_X143Y124_AQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D3 = CLBLM_L_X90Y123_SLICE_X142Y123_B5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D4 = CLBLM_L_X90Y125_SLICE_X142Y125_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_D6 = CLBLM_L_X90Y128_SLICE_X143Y128_BQ;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A1 = CLBLM_L_X90Y128_SLICE_X142Y128_CO6;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A4 = CLBLM_L_X90Y124_SLICE_X142Y124_BO6;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A5 = CLBLM_L_X90Y123_SLICE_X142Y123_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A2 = CLBLL_L_X100Y120_SLICE_X157Y120_A5Q;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A3 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_AX = CLBLM_L_X90Y124_SLICE_X142Y124_BO5;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_A4 = CLBLM_L_X98Y117_SLICE_X155Y117_A5Q;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C5 = CLBLL_L_X102Y125_SLICE_X160Y125_B5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B1 = CLBLM_L_X90Y124_SLICE_X142Y124_AQ;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B2 = CLBLM_L_X90Y124_SLICE_X142Y124_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B4 = CLBLM_L_X90Y124_SLICE_X142Y124_CQ;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B3 = CLBLL_L_X100Y119_SLICE_X157Y119_C5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B5 = CLBLM_L_X90Y124_SLICE_X142Y124_C5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_B6 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C2 = CLBLM_L_X90Y124_SLICE_X142Y124_CQ;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C3 = CLBLM_L_X90Y124_SLICE_X142Y124_AQ;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C5 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C4 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_C6 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B5 = CLBLL_L_X100Y120_SLICE_X156Y120_AQ;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_B6 = 1'b1;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C1 = CLBLL_L_X100Y120_SLICE_X156Y120_AQ;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C3 = CLBLL_L_X102Y120_SLICE_X160Y120_B5Q;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C4 = CLBLL_L_X100Y120_SLICE_X157Y120_BQ;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C5 = CLBLL_L_X100Y119_SLICE_X157Y119_C5Q;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_C6 = CLBLL_L_X100Y119_SLICE_X156Y119_BQ;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D2 = CLBLM_L_X90Y124_SLICE_X142Y124_CQ;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D3 = CLBLM_L_X90Y124_SLICE_X142Y124_AQ;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D5 = CLBLM_L_X92Y122_SLICE_X145Y122_C5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D4 = CLBLM_L_X90Y124_SLICE_X142Y124_A5Q;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D1 = CLBLM_L_X98Y120_SLICE_X155Y120_DO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D4 = CLBLM_R_X101Y125_SLICE_X158Y125_CO6;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D5 = CLBLM_R_X97Y120_SLICE_X153Y120_A5Q;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_D6 = CLBLL_L_X100Y122_SLICE_X157Y122_BQ;
  assign CLBLL_L_X100Y120_SLICE_X157Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D5 = CLBLL_L_X102Y125_SLICE_X160Y125_B5Q;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_A4 = CLBLM_L_X90Y118_SLICE_X142Y118_AQ;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A2 = CLBLM_R_X101Y117_SLICE_X159Y117_AQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A4 = CLBLM_R_X101Y115_SLICE_X158Y115_CO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_AX = CLBLM_L_X98Y134_SLICE_X154Y134_BO5;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B3 = CLBLM_R_X101Y113_SLICE_X159Y113_AQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B4 = CLBLM_R_X101Y116_SLICE_X159Y116_DO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B1 = CLBLM_L_X98Y134_SLICE_X154Y134_CQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B2 = CLBLM_L_X98Y134_SLICE_X154Y134_A5Q;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C2 = CLBLM_R_X101Y116_SLICE_X159Y116_CQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C4 = CLBLL_L_X100Y116_SLICE_X157Y116_BQ;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B3 = CLBLM_L_X98Y134_SLICE_X154Y134_AQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B5 = CLBLM_L_X98Y134_SLICE_X154Y134_C5Q;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D1 = CLBLM_R_X101Y116_SLICE_X159Y116_C5Q;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D2 = CLBLL_L_X100Y116_SLICE_X157Y116_BQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D4 = CLBLM_R_X101Y118_SLICE_X159Y118_A5Q;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_B6 = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D5 = CLBLM_R_X101Y116_SLICE_X159Y116_CQ;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_B5 = CLBLM_L_X90Y117_SLICE_X142Y117_AQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A2 = CLBLL_L_X100Y115_SLICE_X156Y115_CQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A3 = CLBLL_L_X100Y116_SLICE_X156Y116_B5Q;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B2 = CLBLM_R_X101Y116_SLICE_X158Y116_BQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B3 = CLBLM_R_X101Y116_SLICE_X158Y116_AQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C1 = CLBLM_R_X101Y113_SLICE_X159Y113_AQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C2 = CLBLM_R_X101Y114_SLICE_X158Y114_B5Q;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C3 = CLBLM_R_X101Y116_SLICE_X159Y116_DO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C6 = CLBLL_L_X100Y116_SLICE_X157Y116_DO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C3 = CLBLM_L_X98Y134_SLICE_X154Y134_AQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D2 = CLBLM_R_X101Y116_SLICE_X158Y116_AQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D3 = CLBLM_R_X101Y116_SLICE_X158Y116_BQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D4 = CLBLL_L_X100Y115_SLICE_X156Y115_CQ;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C5 = CLBLM_L_X98Y134_SLICE_X154Y134_CQ;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D5 = CLBLM_R_X101Y116_SLICE_X158Y116_B5Q;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_C6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y103_IOB_X1Y104_O = 1'b0;
  assign RIOB33_X105Y103_IOB_X1Y103_O = 1'b0;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y103_IOB_X1Y104_T = 1'b1;
  assign RIOB33_X105Y103_IOB_X1Y103_T = 1'b1;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A3 = CLBLL_L_X100Y120_SLICE_X157Y120_AQ;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A5 = CLBLL_L_X100Y121_SLICE_X156Y121_A5Q;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B3 = CLBLL_L_X100Y121_SLICE_X157Y121_AO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B5 = CLBLM_R_X93Y121_SLICE_X146Y121_DO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D1 = CLBLM_L_X90Y119_SLICE_X143Y119_AQ;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B6 = CLBLL_L_X100Y121_SLICE_X156Y121_A5Q;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C1 = CLBLM_R_X101Y121_SLICE_X159Y121_C5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A1 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A2 = CLBLM_L_X90Y125_SLICE_X143Y125_A5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A4 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A5 = CLBLM_L_X90Y123_SLICE_X142Y123_AQ;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_A6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D5 = CLBLM_L_X98Y134_SLICE_X154Y134_CQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A6 = CLBLL_L_X102Y123_SLICE_X161Y123_CO6;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_D2 = CLBLM_R_X95Y118_SLICE_X150Y118_C5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B1 = CLBLM_L_X90Y116_SLICE_X143Y116_B5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B2 = CLBLM_L_X90Y124_SLICE_X143Y124_AQ;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B4 = CLBLM_R_X89Y125_SLICE_X140Y125_B5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B5 = CLBLM_L_X90Y128_SLICE_X143Y128_DQ;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_B6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D1 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C2 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C3 = CLBLM_L_X92Y131_SLICE_X144Y131_C5Q;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C4 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C5 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_C6 = CLBLM_R_X89Y124_SLICE_X140Y124_BQ;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D2 = CLBLM_L_X90Y125_SLICE_X143Y125_CQ;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D3 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B4 = CLBLL_L_X102Y125_SLICE_X160Y125_B5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D5 = CLBLM_L_X90Y116_SLICE_X143Y116_B5Q;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_D6 = CLBLM_L_X90Y122_SLICE_X143Y122_A5Q;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B5 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X143Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y119_SLICE_X142Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A1 = CLBLL_L_X100Y121_SLICE_X157Y121_CQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B6 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A4 = CLBLM_L_X90Y124_SLICE_X143Y124_BQ;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A5 = CLBLM_R_X89Y125_SLICE_X140Y125_BQ;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A3 = CLBLL_L_X100Y121_SLICE_X157Y121_AQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A4 = CLBLL_L_X100Y121_SLICE_X156Y121_BQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A5 = CLBLM_L_X98Y121_SLICE_X155Y121_C5Q;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B3 = CLBLM_L_X90Y125_SLICE_X142Y125_AQ;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B4 = CLBLM_R_X89Y125_SLICE_X141Y125_C5Q;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B5 = CLBLM_R_X89Y125_SLICE_X140Y125_BQ;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B6 = CLBLM_R_X89Y125_SLICE_X140Y125_B5Q;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B3 = CLBLM_R_X93Y121_SLICE_X147Y121_DO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B4 = CLBLL_L_X102Y121_SLICE_X160Y121_AO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B5 = CLBLL_L_X100Y120_SLICE_X157Y120_AQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C2 = CLBLM_R_X101Y120_SLICE_X158Y120_CQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C5 = CLBLL_L_X100Y121_SLICE_X156Y121_BQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C6 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C1 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C3 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C4 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D1 = CLBLM_L_X98Y121_SLICE_X155Y121_C5Q;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D2 = CLBLL_L_X100Y121_SLICE_X157Y121_CQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D4 = CLBLL_L_X102Y120_SLICE_X160Y120_DQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D5 = CLBLL_L_X100Y121_SLICE_X157Y121_AQ;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D6 = CLBLL_L_X100Y121_SLICE_X156Y121_BQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C4 = CLBLL_L_X102Y125_SLICE_X161Y125_BQ;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C5 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D4 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D5 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C6 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C4 = CLBLM_R_X97Y118_SLICE_X152Y118_A5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C5 = CLBLM_R_X97Y117_SLICE_X152Y117_B5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A3 = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A4 = CLBLL_L_X102Y117_SLICE_X161Y117_AQ;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A6 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B2 = CLBLL_L_X102Y117_SLICE_X160Y117_AQ;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B3 = CLBLM_R_X101Y118_SLICE_X158Y118_B5Q;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C3 = CLBLM_R_X101Y114_SLICE_X158Y114_B5Q;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C4 = CLBLM_R_X101Y118_SLICE_X159Y118_B5Q;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A6 = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_D1 = 1'b0;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_T1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D6 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A1 = CLBLL_L_X100Y118_SLICE_X157Y118_C5Q;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A2 = CLBLM_R_X101Y117_SLICE_X159Y117_B5Q;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A5 = CLBLM_R_X101Y117_SLICE_X159Y117_CQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B1 = CLBLM_R_X101Y115_SLICE_X158Y115_B5Q;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B2 = CLBLM_R_X101Y117_SLICE_X158Y117_BQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B3 = CLBLM_R_X101Y117_SLICE_X158Y117_AQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B4 = CLBLL_L_X102Y116_SLICE_X161Y116_A5Q;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B6 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C1 = CLBLM_R_X101Y117_SLICE_X159Y117_AQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C2 = CLBLL_L_X100Y118_SLICE_X156Y118_CO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C3 = CLBLM_R_X101Y117_SLICE_X158Y117_BQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C6 = CLBLM_R_X101Y115_SLICE_X158Y115_CO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y105_IOB_X1Y106_O = 1'b0;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y105_IOB_X1Y105_O = 1'b0;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D1 = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D2 = CLBLM_R_X101Y117_SLICE_X158Y117_AQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D3 = CLBLM_R_X97Y117_SLICE_X152Y117_DO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D5 = CLBLL_L_X102Y117_SLICE_X161Y117_AQ;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOB33_X105Y105_IOB_X1Y106_T = 1'b1;
  assign RIOB33_X105Y105_IOB_X1Y105_T = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C1 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C2 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D3 = CLBLM_R_X89Y122_SLICE_X141Y122_BQ;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C5 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D4 = CLBLM_R_X89Y122_SLICE_X141Y122_DQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = 1'b0;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D5 = CLBLM_R_X89Y122_SLICE_X141Y122_B5Q;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_C5 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A2 = CLBLL_L_X100Y122_SLICE_X156Y122_A5Q;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D6 = CLBLM_R_X89Y120_SLICE_X141Y120_CQ;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A3 = CLBLM_L_X98Y122_SLICE_X155Y122_AQ;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A4 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A5 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_A6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_R_X103Y124_SLICE_X162Y124_CO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B2 = CLBLL_L_X100Y121_SLICE_X156Y121_CQ;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B3 = CLBLM_R_X101Y122_SLICE_X159Y122_DO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B4 = CLBLM_R_X101Y121_SLICE_X158Y121_CO6;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B5 = CLBLL_L_X100Y122_SLICE_X156Y122_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = 1'b0;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C1 = CLBLM_L_X98Y122_SLICE_X155Y122_AQ;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C4 = CLBLM_R_X101Y122_SLICE_X158Y122_DO6;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C5 = CLBLM_R_X97Y121_SLICE_X152Y121_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_C6 = CLBLM_R_X97Y122_SLICE_X153Y122_DO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A1 = CLBLM_L_X90Y131_SLICE_X142Y131_DO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A4 = CLBLM_L_X90Y126_SLICE_X143Y126_BO6;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A5 = CLBLM_L_X90Y125_SLICE_X143Y125_A5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_AX = CLBLM_L_X90Y126_SLICE_X143Y126_BO5;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B1 = CLBLM_L_X90Y126_SLICE_X143Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B2 = CLBLM_L_X90Y126_SLICE_X143Y126_A5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D1 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D2 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D3 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D4 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D5 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_D6 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X156Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B4 = CLBLM_L_X90Y126_SLICE_X143Y126_CQ;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B5 = CLBLM_L_X90Y126_SLICE_X143Y126_C5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_B6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C2 = CLBLM_L_X90Y126_SLICE_X143Y126_CQ;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C3 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C4 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C5 = CLBLM_L_X90Y126_SLICE_X143Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_C6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y119_SLICE_X146Y119_D1 = CLBLM_R_X93Y119_SLICE_X146Y119_C5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D1 = CLBLM_L_X90Y126_SLICE_X143Y126_C5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D2 = CLBLM_L_X92Y124_SLICE_X145Y124_A5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D4 = CLBLM_L_X90Y126_SLICE_X143Y126_A5Q;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D5 = CLBLM_L_X90Y126_SLICE_X143Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_D6 = CLBLM_L_X90Y126_SLICE_X143Y126_CQ;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_D1 = 1'b0;
  assign CLBLM_L_X90Y126_SLICE_X143Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A1 = CLBLM_R_X101Y122_SLICE_X159Y122_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A2 = CLBLL_L_X100Y122_SLICE_X156Y122_BO6;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A4 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A5 = CLBLL_L_X100Y123_SLICE_X156Y123_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_A6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A4 = CLBLM_R_X89Y126_SLICE_X140Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A5 = CLBLM_L_X90Y126_SLICE_X142Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A1 = CLBLM_L_X90Y126_SLICE_X142Y126_B5Q;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A2 = CLBLM_L_X90Y126_SLICE_X142Y126_BQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B2 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B3 = CLBLL_L_X100Y122_SLICE_X157Y122_CQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B4 = CLBLM_R_X89Y126_SLICE_X140Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B1 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B2 = CLBLM_L_X90Y126_SLICE_X142Y126_BQ;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B4 = CLBLL_L_X100Y122_SLICE_X157Y122_B5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_B5 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_B5 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C1 = CLBLM_R_X101Y122_SLICE_X158Y122_AQ;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C2 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C4 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C5 = CLBLL_L_X100Y122_SLICE_X157Y122_C5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_C6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C4 = CLBLM_L_X92Y124_SLICE_X144Y124_A5Q;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C5 = CLBLM_L_X90Y123_SLICE_X142Y123_C5Q;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C6 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_C2 = CLBLM_L_X90Y126_SLICE_X143Y126_A5Q;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D1 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D2 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D3 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D4 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D5 = 1'b1;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_D6 = 1'b1;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y122_SLICE_X157Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D1 = CLBLM_L_X90Y126_SLICE_X142Y126_BQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D2 = CLBLM_L_X90Y126_SLICE_X142Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D4 = CLBLM_L_X92Y123_SLICE_X144Y123_DQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D5 = CLBLM_L_X90Y126_SLICE_X142Y126_B5Q;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_D6 = CLBLM_R_X89Y126_SLICE_X140Y126_AQ;
  assign CLBLM_L_X90Y126_SLICE_X142Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B6 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C5 = CLBLM_L_X94Y124_SLICE_X149Y124_AQ;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C3 = CLBLM_R_X89Y121_SLICE_X140Y121_AQ;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C4 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A2 = CLBLL_L_X100Y118_SLICE_X157Y118_AQ;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A3 = CLBLM_R_X101Y116_SLICE_X159Y116_C5Q;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A4 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B2 = CLBLM_R_X101Y118_SLICE_X159Y118_BQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B3 = CLBLM_R_X101Y118_SLICE_X159Y118_AQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B4 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C2 = CLBLM_R_X101Y118_SLICE_X159Y118_CQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C3 = CLBLM_L_X98Y117_SLICE_X155Y117_DO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C5 = CLBLM_R_X101Y118_SLICE_X159Y118_DO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C6 = CLBLM_R_X101Y117_SLICE_X159Y117_CQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_CX = CLBLM_R_X101Y116_SLICE_X159Y116_BO5;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D2 = CLBLM_R_X101Y118_SLICE_X159Y118_AQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D3 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D4 = CLBLM_R_X101Y118_SLICE_X159Y118_BQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D5 = CLBLM_R_X101Y118_SLICE_X159Y118_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D6 = CLBLL_L_X100Y118_SLICE_X157Y118_AQ;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A2 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A3 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A4 = CLBLM_R_X101Y117_SLICE_X158Y117_DO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A5 = CLBLL_L_X100Y120_SLICE_X157Y120_DO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A6 = 1'b1;
  assign RIOB33_X105Y107_IOB_X1Y107_O = 1'b0;
  assign RIOB33_X105Y107_IOB_X1Y108_O = 1'b0;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B2 = CLBLM_R_X101Y118_SLICE_X158Y118_BQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B3 = CLBLM_R_X101Y118_SLICE_X158Y118_AQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B4 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B6 = 1'b1;
  assign RIOB33_X105Y107_IOB_X1Y107_T = 1'b1;
  assign RIOB33_X105Y107_IOB_X1Y108_T = 1'b1;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_D1 = 1'b0;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C1 = CLBLL_L_X102Y117_SLICE_X160Y117_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C2 = CLBLM_R_X101Y119_SLICE_X158Y119_CQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C4 = CLBLM_R_X101Y117_SLICE_X159Y117_CQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D5 = CLBLM_R_X89Y120_SLICE_X140Y120_CQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_T1 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D2 = CLBLM_R_X101Y118_SLICE_X158Y118_AQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D3 = CLBLM_R_X101Y117_SLICE_X159Y117_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D4 = CLBLM_R_X101Y118_SLICE_X158Y118_BQ;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D5 = CLBLM_R_X101Y118_SLICE_X158Y118_B5Q;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A2 = CLBLM_R_X101Y123_SLICE_X158Y123_B5Q;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A3 = CLBLL_L_X100Y122_SLICE_X156Y122_CO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A4 = CLBLL_L_X100Y123_SLICE_X156Y123_B5Q;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B2 = CLBLM_L_X98Y125_SLICE_X154Y125_A5Q;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B3 = CLBLM_L_X98Y122_SLICE_X155Y122_CO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B4 = CLBLM_R_X101Y123_SLICE_X158Y123_A5Q;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A2 = CLBLL_L_X100Y123_SLICE_X157Y123_A5Q;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A3 = CLBLL_L_X100Y122_SLICE_X157Y122_BQ;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C6 = 1'b1;
  assign LIOB33_X0Y239_IOB_X0Y240_T = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A3 = CLBLM_R_X101Y120_SLICE_X159Y120_B5Q;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A4 = CLBLM_R_X101Y119_SLICE_X158Y119_BQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B2 = CLBLM_R_X101Y119_SLICE_X159Y119_BQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B3 = CLBLM_R_X101Y119_SLICE_X159Y119_AQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B6 = 1'b1;
  assign RIOB33_X105Y109_IOB_X1Y109_O = CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C1 = CLBLL_L_X102Y117_SLICE_X161Y117_CQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C3 = CLBLM_R_X101Y119_SLICE_X159Y119_BQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C4 = CLBLM_R_X101Y119_SLICE_X159Y119_AQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C5 = CLBLM_R_X101Y119_SLICE_X159Y119_B5Q;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C6 = CLBLM_R_X101Y119_SLICE_X158Y119_BQ;
  assign RIOB33_X105Y109_IOB_X1Y110_O = CLBLM_R_X101Y113_SLICE_X159Y113_AO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D1 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D3 = CLBLM_R_X101Y119_SLICE_X159Y119_BQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D4 = CLBLM_R_X101Y119_SLICE_X159Y119_AQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D5 = CLBLM_R_X101Y119_SLICE_X159Y119_B5Q;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D6 = CLBLM_R_X101Y119_SLICE_X158Y119_BQ;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A3 = CLBLL_L_X100Y119_SLICE_X157Y119_CQ;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A5 = CLBLM_R_X101Y120_SLICE_X158Y120_AQ;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B2 = CLBLM_R_X101Y119_SLICE_X159Y119_DO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B3 = CLBLL_L_X102Y117_SLICE_X161Y117_CQ;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B6 = CLBLM_L_X98Y119_SLICE_X154Y119_DO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C1 = CLBLM_R_X101Y123_SLICE_X159Y123_C5Q;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C2 = CLBLM_R_X101Y119_SLICE_X159Y119_A5Q;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D1 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D3 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = 1'b0;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A2 = CLBLL_L_X100Y125_SLICE_X157Y125_DQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A3 = CLBLL_L_X100Y124_SLICE_X156Y124_B5Q;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A4 = CLBLL_L_X100Y124_SLICE_X156Y124_AQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A5 = CLBLL_L_X100Y124_SLICE_X156Y124_BQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_A6 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B2 = CLBLL_L_X100Y125_SLICE_X157Y125_DQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B3 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B4 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B5 = CLBLL_L_X100Y124_SLICE_X156Y124_BQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_B6 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C1 = CLBLL_L_X100Y124_SLICE_X156Y124_BQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C3 = CLBLM_L_X98Y125_SLICE_X154Y125_D5Q;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C4 = CLBLL_L_X100Y125_SLICE_X157Y125_DQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C5 = CLBLL_L_X100Y124_SLICE_X156Y124_B5Q;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_C6 = CLBLL_L_X100Y124_SLICE_X156Y124_AQ;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y55_IOB_X0Y56_O = 1'b0;
  assign LIOB33_X0Y55_IOB_X0Y55_O = 1'b0;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D1 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A1 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A2 = CLBLM_L_X90Y128_SLICE_X143Y128_A5Q;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D2 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D3 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D4 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D5 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_D6 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X156Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B1 = CLBLM_L_X90Y124_SLICE_X143Y124_AO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B2 = CLBLM_L_X92Y128_SLICE_X145Y128_DO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A5 = CLBLM_R_X89Y127_SLICE_X141Y127_AQ;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B6 = CLBLM_L_X90Y128_SLICE_X143Y128_A5Q;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C2 = CLBLM_L_X90Y128_SLICE_X142Y128_AO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C3 = CLBLM_R_X89Y127_SLICE_X141Y127_AQ;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C4 = CLBLM_L_X92Y129_SLICE_X145Y129_DO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A2 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A3 = CLBLL_L_X100Y124_SLICE_X157Y124_AQ;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A4 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A5 = CLBLL_L_X100Y125_SLICE_X157Y125_AQ;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D1 = CLBLM_L_X90Y128_SLICE_X142Y128_AQ;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D2 = CLBLM_L_X90Y125_SLICE_X143Y125_B5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_A6 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D3 = CLBLM_L_X90Y129_SLICE_X142Y129_A5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D4 = CLBLM_L_X92Y126_SLICE_X145Y126_C5Q;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B4 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B5 = CLBLL_L_X100Y124_SLICE_X157Y124_A5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B6 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B2 = CLBLL_L_X100Y125_SLICE_X157Y125_C5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_B3 = CLBLM_L_X98Y124_SLICE_X154Y124_CO6;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A1 = CLBLM_L_X90Y128_SLICE_X142Y128_B5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C2 = CLBLL_L_X100Y123_SLICE_X157Y123_A5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C3 = CLBLM_L_X98Y124_SLICE_X154Y124_DO6;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A2 = CLBLM_L_X90Y128_SLICE_X142Y128_AQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A4 = CLBLM_R_X89Y128_SLICE_X141Y128_AQ;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C5 = CLBLL_L_X100Y124_SLICE_X157Y124_DO6;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B2 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B4 = CLBLM_R_X89Y128_SLICE_X141Y128_AQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B5 = CLBLM_L_X90Y129_SLICE_X142Y129_AQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B6 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D1 = CLBLL_L_X100Y125_SLICE_X157Y125_AQ;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D2 = CLBLL_L_X100Y126_SLICE_X157Y126_CQ;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D4 = CLBLL_L_X100Y124_SLICE_X157Y124_A5Q;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D5 = 1'b1;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_D6 = CLBLL_L_X100Y124_SLICE_X157Y124_AQ;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C3 = CLBLM_L_X90Y128_SLICE_X142Y128_BQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C4 = CLBLM_L_X90Y129_SLICE_X142Y129_C5Q;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C5 = CLBLM_L_X90Y129_SLICE_X142Y129_A5Q;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C6 = CLBLM_L_X90Y123_SLICE_X142Y123_C5Q;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D1 = CLBLM_L_X90Y123_SLICE_X142Y123_CQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D4 = CLBLM_L_X90Y128_SLICE_X143Y128_CQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D5 = CLBLM_L_X90Y128_SLICE_X142Y128_B5Q;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D6 = CLBLM_R_X89Y128_SLICE_X141Y128_AQ;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_D2 = CLBLM_L_X90Y128_SLICE_X142Y128_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X103Y124_SLICE_X163Y124_CO6;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = 1'b0;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLL_L_X102Y124_SLICE_X161Y124_CO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_D1 = 1'b0;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLM_R_X103Y121_SLICE_X162Y121_CO6;
  assign RIOB33_X105Y111_IOB_X1Y111_O = CLBLM_R_X101Y113_SLICE_X159Y113_BO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A1 = CLBLM_R_X101Y120_SLICE_X159Y120_DO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A2 = CLBLL_L_X102Y122_SLICE_X160Y122_BQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A4 = CLBLM_L_X98Y120_SLICE_X155Y120_CO6;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = 1'b0;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B2 = CLBLM_R_X101Y120_SLICE_X159Y120_BQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B3 = CLBLM_R_X101Y120_SLICE_X159Y120_AQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B4 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B5 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_B6 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C1 = CLBLM_R_X101Y119_SLICE_X159Y119_A5Q;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C2 = CLBLM_R_X101Y120_SLICE_X159Y120_AQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C3 = CLBLM_R_X101Y120_SLICE_X159Y120_BQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C5 = CLBLM_R_X101Y120_SLICE_X159Y120_B5Q;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_C6 = CLBLL_L_X102Y122_SLICE_X160Y122_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = 1'b0;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D1 = CLBLM_R_X101Y120_SLICE_X159Y120_BQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D2 = CLBLM_R_X101Y120_SLICE_X159Y120_AQ;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D3 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D5 = CLBLM_R_X101Y120_SLICE_X159Y120_B5Q;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_D6 = CLBLM_R_X101Y119_SLICE_X159Y119_A5Q;
  assign CLBLM_R_X101Y120_SLICE_X159Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A3 = CLBLL_L_X100Y120_SLICE_X157Y120_A5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A4 = CLBLM_R_X101Y120_SLICE_X158Y120_BO6;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A5 = CLBLM_L_X94Y121_SLICE_X148Y121_DO6;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_AX = CLBLM_R_X101Y120_SLICE_X158Y120_BO5;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B2 = CLBLM_R_X101Y120_SLICE_X158Y120_A5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B3 = CLBLM_R_X101Y119_SLICE_X158Y119_AQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B4 = CLBLM_R_X101Y120_SLICE_X158Y120_AQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B5 = CLBLM_R_X101Y120_SLICE_X158Y120_C5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_B6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A4 = CLBLM_L_X90Y116_SLICE_X143Y116_B5Q;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D4 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C1 = CLBLM_R_X101Y119_SLICE_X158Y119_AQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C2 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D5 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C4 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C5 = CLBLL_L_X100Y121_SLICE_X157Y121_BQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_C6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_A6 = 1'b1;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D1 = CLBLM_R_X101Y120_SLICE_X158Y120_C5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D3 = CLBLM_R_X101Y120_SLICE_X158Y120_AQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D4 = CLBLM_R_X101Y120_SLICE_X158Y120_A5Q;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D5 = CLBLM_R_X101Y119_SLICE_X158Y119_AQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_D6 = CLBLL_L_X102Y120_SLICE_X160Y120_CQ;
  assign CLBLM_R_X101Y120_SLICE_X158Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B4 = CLBLM_L_X90Y119_SLICE_X143Y119_AO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A1 = CLBLL_L_X100Y125_SLICE_X156Y125_DO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A3 = CLBLL_L_X100Y126_SLICE_X157Y126_A5Q;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A5 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_A6 = CLBLL_L_X100Y125_SLICE_X156Y125_CO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_B6 = CLBLM_L_X94Y123_SLICE_X148Y123_DO6;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B2 = CLBLL_L_X100Y125_SLICE_X156Y125_BQ;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B3 = CLBLL_L_X100Y125_SLICE_X156Y125_AQ;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B4 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B5 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_B6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C2 = CLBLL_L_X100Y125_SLICE_X156Y125_AQ;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C3 = CLBLL_L_X100Y125_SLICE_X156Y125_BQ;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C4 = CLBLL_L_X100Y126_SLICE_X156Y126_A5Q;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C5 = CLBLL_L_X100Y125_SLICE_X156Y125_B5Q;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_C6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D2 = CLBLM_L_X98Y125_SLICE_X154Y125_C5Q;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D5 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C3 = CLBLM_L_X90Y120_SLICE_X143Y120_BQ;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A1 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A4 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X156Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C4 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_C5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A2 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_A3 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B2 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B4 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B1 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B6 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B3 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_B5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C1 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C2 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C3 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C4 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_C6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A2 = CLBLL_L_X100Y126_SLICE_X157Y126_CQ;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A3 = CLBLM_R_X101Y125_SLICE_X158Y125_B5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A4 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D1 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D2 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D3 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D4 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X143Y129_D6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_A6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B5 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B2 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B3 = CLBLM_L_X98Y126_SLICE_X154Y126_AQ;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_B4 = CLBLL_L_X100Y125_SLICE_X157Y125_B5Q;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A1 = CLBLM_R_X93Y131_SLICE_X146Y131_DO6;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A2 = CLBLM_L_X90Y128_SLICE_X143Y128_AQ;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C5 = CLBLM_R_X103Y126_SLICE_X163Y126_A5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C6 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A4 = CLBLM_L_X90Y129_SLICE_X142Y129_BO6;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_AX = CLBLM_L_X90Y129_SLICE_X142Y129_BO5;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C2 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C3 = CLBLL_L_X100Y125_SLICE_X157Y125_A5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B1 = CLBLM_L_X90Y129_SLICE_X142Y129_AQ;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B2 = CLBLM_L_X90Y129_SLICE_X142Y129_A5Q;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B4 = CLBLM_L_X90Y128_SLICE_X142Y128_BQ;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B5 = CLBLM_L_X90Y129_SLICE_X142Y129_C5Q;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_B6 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C2 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C4 = CLBLM_L_X90Y128_SLICE_X142Y128_BQ;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D2 = CLBLL_L_X100Y124_SLICE_X156Y124_AO6;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D3 = CLBLL_L_X102Y125_SLICE_X160Y125_DO6;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D5 = CLBLL_L_X100Y125_SLICE_X157Y125_B5Q;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D4 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D1 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D2 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D3 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D6 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D5 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D4 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_D6 = 1'b1;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y59_IOB_X0Y60_O = 1'b0;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A2 = CLBLM_R_X101Y121_SLICE_X158Y121_BO6;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A3 = CLBLM_R_X101Y122_SLICE_X159Y122_B5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A4 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A5 = CLBLL_L_X100Y122_SLICE_X157Y122_A5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_A6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D3 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D4 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B2 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B3 = CLBLM_R_X101Y121_SLICE_X159Y121_AQ;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B4 = CLBLM_R_X101Y121_SLICE_X158Y121_A5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B5 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D5 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_B6 = 1'b1;
  assign LIOB33_X0Y59_IOB_X0Y59_O = 1'b0;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D6 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C2 = CLBLM_R_X101Y121_SLICE_X159Y121_CQ;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C4 = CLBLM_R_X101Y121_SLICE_X159Y121_BQ;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C5 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_C6 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D1 = CLBLM_R_X101Y121_SLICE_X159Y121_C5Q;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D2 = CLBLM_R_X101Y121_SLICE_X159Y121_CQ;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D4 = CLBLM_R_X101Y121_SLICE_X159Y121_BQ;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D5 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_D6 = CLBLM_R_X101Y121_SLICE_X159Y121_AQ;
  assign CLBLM_R_X101Y121_SLICE_X159Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A2 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A3 = CLBLM_R_X101Y121_SLICE_X158Y121_AQ;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A4 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A5 = CLBLL_L_X100Y122_SLICE_X157Y122_AQ;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_A6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B4 = CLBLM_R_X89Y121_SLICE_X140Y121_CQ;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B1 = CLBLL_L_X100Y122_SLICE_X156Y122_AQ;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B2 = CLBLM_R_X101Y121_SLICE_X159Y121_DO6;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B3 = CLBLM_R_X103Y121_SLICE_X163Y121_DO6;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B4 = CLBLL_L_X100Y121_SLICE_X156Y121_C5Q;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C1 = CLBLL_L_X100Y122_SLICE_X157Y122_AQ;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C2 = CLBLM_R_X101Y121_SLICE_X158Y121_AQ;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C3 = CLBLM_R_X101Y121_SLICE_X159Y121_B5Q;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C4 = CLBLM_R_X101Y121_SLICE_X158Y121_A5Q;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C5 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D1 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D2 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D3 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D4 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D5 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_D6 = 1'b1;
  assign CLBLM_R_X101Y121_SLICE_X158Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A4 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A1 = CLBLL_L_X100Y125_SLICE_X156Y125_B5Q;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A2 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A3 = CLBLL_L_X100Y126_SLICE_X157Y126_BQ;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A5 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_A6 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B1 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B2 = CLBLL_L_X100Y126_SLICE_X156Y126_BQ;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B3 = CLBLL_L_X100Y126_SLICE_X156Y126_AQ;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B5 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_B6 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C2 = CLBLL_L_X100Y126_SLICE_X156Y126_AQ;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C3 = CLBLL_L_X100Y126_SLICE_X156Y126_BQ;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C4 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C5 = CLBLL_L_X100Y126_SLICE_X156Y126_B5Q;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_C6 = CLBLL_L_X100Y126_SLICE_X157Y126_BQ;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_A6 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D3 = CLBLM_L_X98Y126_SLICE_X154Y126_B5Q;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D5 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y126_SLICE_X156Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A1 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A2 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A3 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A4 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A5 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_A6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D2 = CLBLM_R_X89Y120_SLICE_X141Y120_AQ;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B1 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B2 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B3 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B5 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B2 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B6 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_B4 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C1 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C2 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C3 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C4 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C5 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A2 = CLBLL_L_X100Y126_SLICE_X157Y126_A5Q;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A3 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_C6 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A5 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A6 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B5 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B1 = CLBLL_L_X100Y126_SLICE_X157Y126_AQ;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_A4 = CLBLM_R_X101Y126_SLICE_X158Y126_AQ;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B3 = CLBLL_L_X100Y126_SLICE_X156Y126_CO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B6 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D1 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D2 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D3 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D4 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C2 = CLBLM_R_X101Y126_SLICE_X158Y126_BO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C4 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D6 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A2 = CLBLM_L_X90Y130_SLICE_X142Y130_A5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A3 = CLBLM_L_X90Y128_SLICE_X143Y128_AQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A4 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A5 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_A6 = 1'b1;
  assign CLBLM_L_X90Y120_SLICE_X142Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B2 = CLBLM_L_X90Y130_SLICE_X142Y130_A5Q;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B6 = CLBLM_L_X90Y130_SLICE_X142Y130_CO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C1 = CLBLL_L_X102Y128_SLICE_X161Y128_AQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_B3 = CLBLM_L_X92Y131_SLICE_X144Y131_DO6;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_BX = CLBLM_L_X90Y130_SLICE_X142Y130_CO5;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D2 = CLBLM_L_X98Y127_SLICE_X155Y127_CO6;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C2 = CLBLL_L_X102Y126_SLICE_X160Y126_C5Q;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D4 = CLBLM_L_X98Y125_SLICE_X154Y125_A5Q;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D6 = CLBLL_L_X100Y125_SLICE_X157Y125_BQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C1 = CLBLM_L_X90Y131_SLICE_X142Y131_C5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C2 = CLBLM_L_X90Y130_SLICE_X142Y130_B5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C3 = CLBLM_L_X90Y129_SLICE_X142Y129_CQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C4 = CLBLM_L_X90Y130_SLICE_X142Y130_BQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_C6 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C5 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C6 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D1 = CLBLM_L_X90Y131_SLICE_X142Y131_C5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D2 = CLBLM_L_X90Y126_SLICE_X142Y126_CQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D3 = CLBLM_L_X90Y129_SLICE_X142Y129_CQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D4 = CLBLM_L_X90Y130_SLICE_X142Y130_BQ;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D5 = CLBLM_L_X90Y130_SLICE_X142Y130_B5Q;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y130_SLICE_X142Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C4 = CLBLM_R_X97Y118_SLICE_X153Y118_AQ;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C5 = CLBLM_R_X97Y119_SLICE_X152Y119_CQ;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A2 = CLBLL_L_X102Y122_SLICE_X161Y122_CQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A3 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A4 = CLBLM_R_X101Y122_SLICE_X158Y122_B5Q;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A5 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_A6 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B2 = CLBLM_R_X101Y122_SLICE_X159Y122_BQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B3 = CLBLM_R_X101Y122_SLICE_X159Y122_AQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B4 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B5 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_B6 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C1 = CLBLM_R_X101Y122_SLICE_X158Y122_AQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C2 = CLBLM_R_X101Y121_SLICE_X159Y121_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C3 = CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C5 = CLBLM_R_X101Y122_SLICE_X159Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A4 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A5 = CLBLM_R_X101Y135_SLICE_X159Y135_AQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A6 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D2 = CLBLM_R_X101Y122_SLICE_X159Y122_AQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D3 = CLBLM_R_X101Y122_SLICE_X159Y122_BQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D4 = CLBLL_L_X102Y122_SLICE_X161Y122_CQ;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D5 = CLBLM_R_X101Y122_SLICE_X159Y122_B5Q;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_D6 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_BX = CLBLM_R_X89Y122_SLICE_X141Y122_CO5;
  assign CLBLM_R_X101Y122_SLICE_X159Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = 1'b0;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A2 = CLBLM_R_X101Y122_SLICE_X158Y122_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A3 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A4 = CLBLM_R_X101Y124_SLICE_X158Y124_AQ;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A5 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_A6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B2 = CLBLM_R_X101Y122_SLICE_X158Y122_BQ;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B3 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B4 = CLBLL_L_X102Y122_SLICE_X160Y122_CQ;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B5 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_B6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = 1'b0;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C3 = CLBLL_L_X102Y122_SLICE_X161Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C4 = CLBLM_R_X101Y122_SLICE_X158Y122_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C5 = CLBLL_L_X100Y122_SLICE_X157Y122_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_C6 = CLBLM_R_X101Y122_SLICE_X158Y122_DO6;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D2 = CLBLM_R_X101Y122_SLICE_X159Y122_A5Q;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D3 = CLBLM_R_X101Y122_SLICE_X158Y122_BQ;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D4 = 1'b1;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D5 = CLBLM_R_X101Y122_SLICE_X158Y122_B5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_D6 = CLBLL_L_X102Y122_SLICE_X160Y122_CQ;
  assign CLBLM_R_X101Y122_SLICE_X158Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y124_SLICE_X157Y124_C6 = CLBLM_R_X97Y121_SLICE_X153Y121_B5Q;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A1 = CLBLL_L_X100Y127_SLICE_X156Y127_B5Q;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A3 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A4 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A5 = CLBLL_L_X100Y127_SLICE_X157Y127_AQ;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_A6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C1 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_D1 = 1'b0;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C2 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B1 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B3 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B4 = CLBLL_L_X100Y128_SLICE_X156Y128_BQ;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B5 = CLBLL_L_X100Y127_SLICE_X156Y127_BQ;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_B6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_T1 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D2 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C4 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C2 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C3 = CLBLL_L_X100Y127_SLICE_X156Y127_BQ;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C4 = CLBLL_L_X100Y127_SLICE_X156Y127_A5Q;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C5 = CLBLL_L_X100Y127_SLICE_X156Y127_B5Q;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_C6 = CLBLL_L_X100Y128_SLICE_X156Y128_BQ;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = 1'b0;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D1 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D2 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D3 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D4 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D5 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_D6 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X156Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A1 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A2 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A3 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A4 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A5 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_A6 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B1 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B2 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B3 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B4 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B5 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_B6 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A2 = CLBLL_L_X100Y129_SLICE_X157Y129_BO6;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A4 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A5 = CLBLL_L_X100Y128_SLICE_X156Y128_AQ;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_A6 = CLBLL_L_X100Y127_SLICE_X157Y127_CO6;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C1 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C2 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_C3 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B1 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B2 = CLBLL_L_X100Y127_SLICE_X157Y127_BQ;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B3 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B5 = CLBLL_L_X100Y127_SLICE_X156Y127_AQ;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_B6 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D1 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D2 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C1 = CLBLL_L_X100Y127_SLICE_X156Y127_AQ;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C2 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C3 = CLBLL_L_X100Y127_SLICE_X157Y127_BQ;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C4 = CLBLL_L_X100Y127_SLICE_X157Y127_AQ;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C5 = CLBLL_L_X100Y127_SLICE_X157Y127_B5Q;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D3 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D4 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D5 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X143Y131_D6 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A1 = CLBLM_R_X93Y133_SLICE_X146Y133_DO6;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D1 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D2 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D3 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D4 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D5 = 1'b1;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_D6 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_AX = CLBLM_L_X90Y131_SLICE_X142Y131_BO5;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B1 = CLBLM_R_X89Y131_SLICE_X140Y131_A5Q;
  assign CLBLL_L_X100Y127_SLICE_X157Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B2 = CLBLM_L_X90Y131_SLICE_X142Y131_A5Q;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B3 = CLBLM_L_X90Y131_SLICE_X142Y131_AQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B4 = CLBLM_L_X90Y131_SLICE_X142Y131_CQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_B6 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C2 = CLBLM_L_X90Y131_SLICE_X142Y131_AQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C3 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C4 = CLBLM_L_X90Y129_SLICE_X142Y129_CQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C5 = 1'b1;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_C6 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_AX = CLBLM_R_X89Y122_SLICE_X140Y122_BO5;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_D1 = 1'b0;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D1 = CLBLM_L_X90Y126_SLICE_X142Y126_C5Q;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D2 = CLBLM_L_X90Y131_SLICE_X142Y131_CQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D3 = CLBLM_L_X90Y131_SLICE_X142Y131_AQ;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D4 = CLBLM_L_X90Y131_SLICE_X142Y131_A5Q;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D5 = CLBLM_R_X89Y131_SLICE_X140Y131_A5Q;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b0;
  assign CLBLM_L_X90Y131_SLICE_X142Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign RIOI3_X105Y77_ILOGIC_X1Y78_D = RIOB33_X105Y77_IOB_X1Y78_I;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A1 = CLBLL_L_X102Y126_SLICE_X160Y126_AQ;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A5 = CLBLM_R_X101Y123_SLICE_X159Y123_A5Q;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B1 = CLBLL_L_X102Y122_SLICE_X160Y122_DO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B5 = CLBLL_L_X102Y123_SLICE_X161Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B6 = CLBLM_R_X101Y123_SLICE_X159Y123_A5Q;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C1 = CLBLL_L_X102Y124_SLICE_X160Y124_C5Q;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C2 = CLBLL_L_X102Y124_SLICE_X160Y124_D5Q;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C4 = CLBLL_L_X102Y123_SLICE_X160Y123_B5Q;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C5 = CLBLM_R_X101Y123_SLICE_X159Y123_CQ;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A3 = CLBLM_R_X101Y124_SLICE_X158Y124_B5Q;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A4 = CLBLL_L_X102Y123_SLICE_X161Y123_AQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B2 = CLBLM_R_X101Y123_SLICE_X158Y123_BQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B3 = CLBLM_R_X101Y123_SLICE_X158Y123_AQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C3 = CLBLL_L_X102Y122_SLICE_X160Y122_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C4 = CLBLM_R_X101Y124_SLICE_X158Y124_AQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C5 = CLBLL_L_X100Y123_SLICE_X156Y123_A5Q;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C6 = CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D2 = CLBLM_R_X101Y123_SLICE_X158Y123_AQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D3 = CLBLM_R_X101Y123_SLICE_X158Y123_BQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D5 = CLBLM_R_X101Y123_SLICE_X158Y123_B5Q;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D6 = CLBLL_L_X102Y123_SLICE_X161Y123_AQ;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A2 = CLBLL_L_X100Y128_SLICE_X156Y128_A5Q;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A4 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A5 = CLBLL_L_X100Y126_SLICE_X157Y126_AQ;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_A6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B2 = CLBLL_L_X100Y127_SLICE_X156Y127_CO6;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B5 = CLBLL_L_X100Y128_SLICE_X156Y128_A5Q;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_B6 = CLBLL_L_X100Y128_SLICE_X156Y128_CO6;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_B2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_C6 = CLBLM_L_X98Y127_SLICE_X154Y127_B5Q;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C3 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C4 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_C5 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D4 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D5 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_D6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X156Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D3 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D4 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_D5 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A2 = CLBLM_R_X97Y112_SLICE_X153Y112_BQ;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A3 = CLBLM_L_X98Y110_SLICE_X154Y110_AQ;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A4 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A5 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_A6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B1 = CLBLM_L_X98Y111_SLICE_X154Y111_A5Q;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B3 = CLBLM_L_X98Y110_SLICE_X154Y110_AQ;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B4 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B5 = CLBLM_R_X97Y112_SLICE_X153Y112_BQ;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_B6 = CLBLM_L_X98Y110_SLICE_X154Y110_A5Q;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A4 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A5 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_A6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_C2 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B4 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B5 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_B6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D1 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C4 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C5 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_C6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D4 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D5 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_D6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X154Y110_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D1 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D2 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D3 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D4 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D5 = 1'b1;
  assign CLBLL_L_X100Y128_SLICE_X157Y128_D6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = 1'b0;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A3 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A4 = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_D1 = 1'b0;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A2 = CLBLL_L_X102Y126_SLICE_X161Y126_C5Q;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A3 = CLBLM_R_X101Y124_SLICE_X158Y124_CO6;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A4 = CLBLL_L_X102Y126_SLICE_X161Y126_D5Q;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A5 = CLBLM_R_X101Y128_SLICE_X158Y128_A5Q;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_A6 = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_T1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_B6 = 1'b1;
  assign LIOB33_X0Y57_IOB_X0Y57_O = 1'b0;
  assign LIOB33_X0Y57_IOB_X0Y58_O = 1'b0;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_C6 = 1'b1;
  assign CLBLM_L_X98Y110_SLICE_X155Y110_A6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D1 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D2 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_D6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X159Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A2 = CLBLM_R_X101Y124_SLICE_X158Y124_A5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A4 = CLBLL_L_X100Y125_SLICE_X157Y125_BQ;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A5 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_A6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B2 = CLBLM_R_X101Y124_SLICE_X158Y124_BQ;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B3 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B4 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B5 = CLBLM_R_X101Y124_SLICE_X159Y124_AQ;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_B6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C3 = CLBLL_L_X100Y123_SLICE_X156Y123_B5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C4 = CLBLM_R_X101Y124_SLICE_X158Y124_A5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C5 = CLBLM_R_X101Y124_SLICE_X158Y124_DO6;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_C6 = CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  assign LIOB33_X0Y57_IOB_X0Y57_T = 1'b1;
  assign LIOB33_X0Y57_IOB_X0Y58_T = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D2 = CLBLM_R_X101Y123_SLICE_X158Y123_A5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D3 = CLBLM_R_X101Y124_SLICE_X159Y124_AQ;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D4 = CLBLM_R_X101Y124_SLICE_X158Y124_BQ;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D5 = CLBLM_R_X101Y124_SLICE_X158Y124_B5Q;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_D6 = 1'b1;
  assign CLBLM_R_X101Y124_SLICE_X158Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A1 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A3 = CLBLL_L_X100Y130_SLICE_X156Y130_AQ;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A4 = CLBLM_L_X98Y128_SLICE_X154Y128_A5Q;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A5 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_A6 = CLBLM_R_X97Y128_SLICE_X153Y128_A5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A2 = CLBLL_L_X100Y111_SLICE_X156Y111_CO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A3 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B2 = CLBLM_L_X98Y128_SLICE_X154Y128_A5Q;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B4 = CLBLM_R_X101Y129_SLICE_X158Y129_CO6;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B5 = CLBLM_L_X98Y129_SLICE_X155Y129_AQ;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_B6 = CLBLM_L_X98Y128_SLICE_X154Y128_DO6;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A4 = CLBLM_L_X98Y111_SLICE_X155Y111_B5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A5 = CLBLL_L_X100Y111_SLICE_X157Y111_B5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_A6 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C1 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C2 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C3 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C4 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C5 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_C6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B3 = CLBLM_R_X97Y111_SLICE_X152Y111_B5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B4 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_B6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C1 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C2 = CLBLM_L_X98Y111_SLICE_X155Y111_CQ;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D1 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D2 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D3 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D4 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D5 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_D6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y129_SLICE_X156Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D1 = CLBLM_L_X98Y111_SLICE_X155Y111_C5Q;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D2 = CLBLM_L_X98Y111_SLICE_X155Y111_CQ;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D4 = CLBLM_L_X98Y111_SLICE_X155Y111_BQ;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D5 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_D6 = CLBLM_R_X95Y111_SLICE_X150Y111_AQ;
  assign CLBLM_L_X98Y111_SLICE_X155Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A2 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A3 = CLBLM_L_X98Y110_SLICE_X154Y110_A5Q;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A4 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A5 = CLBLM_R_X97Y112_SLICE_X152Y112_AQ;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_A6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = 1'b0;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B2 = CLBLM_L_X98Y111_SLICE_X154Y111_BQ;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B3 = CLBLM_L_X98Y111_SLICE_X154Y111_AQ;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B4 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B5 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_B6 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A2 = CLBLL_L_X100Y129_SLICE_X156Y129_BO6;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A3 = CLBLM_L_X98Y127_SLICE_X155Y127_A5Q;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A4 = CLBLM_R_X101Y130_SLICE_X158Y130_C5Q;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A5 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_A6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C1 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C3 = CLBLM_R_X97Y112_SLICE_X152Y112_AQ;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B2 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B4 = CLBLM_L_X98Y127_SLICE_X155Y127_A5Q;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C4 = CLBLM_L_X98Y111_SLICE_X154Y111_BQ;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C1 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C2 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C3 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C4 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C5 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_C6 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D1 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D2 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D3 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D4 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D5 = 1'b1;
  assign CLBLM_L_X98Y111_SLICE_X154Y111_D6 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D1 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D2 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D3 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D4 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D5 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_D6 = 1'b1;
  assign CLBLL_L_X100Y129_SLICE_X157Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X103Y120_SLICE_X163Y120_CO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLL_L_X102Y118_SLICE_X160Y118_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign LIOB33_X0Y201_IOB_X0Y202_O = 1'b0;
  assign LIOB33_X0Y201_IOB_X0Y201_O = 1'b0;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A1 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A2 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A3 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A4 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_A6 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B1 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B2 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B3 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B4 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_B6 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = 1'b0;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C1 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C2 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C3 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C4 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_C6 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D1 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D2 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D3 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D4 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X159Y125_D6 = 1'b1;
  assign LIOI3_SING_X0Y249_OLOGIC_X0Y249_D1 = 1'b0;
  assign LIOB33_X0Y201_IOB_X0Y202_T = 1'b1;
  assign LIOI3_SING_X0Y249_OLOGIC_X0Y249_T1 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A1 = CLBLM_R_X101Y125_SLICE_X158Y125_DO6;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A3 = CLBLM_R_X101Y126_SLICE_X158Y126_A5Q;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_A6 = CLBLM_R_X101Y125_SLICE_X158Y125_CO6;
  assign LIOB33_X0Y201_IOB_X0Y201_T = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B2 = CLBLM_R_X101Y125_SLICE_X158Y125_BQ;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B3 = CLBLM_R_X101Y125_SLICE_X158Y125_AQ;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B4 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_B6 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C2 = CLBLM_R_X101Y125_SLICE_X158Y125_AQ;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C3 = CLBLL_L_X100Y125_SLICE_X157Y125_A5Q;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C4 = CLBLM_R_X101Y125_SLICE_X158Y125_BQ;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C5 = CLBLM_R_X101Y125_SLICE_X158Y125_B5Q;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_C6 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D5 = 1'b1;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_D6 = CLBLL_L_X100Y125_SLICE_X157Y125_C5Q;
  assign CLBLM_R_X101Y125_SLICE_X158Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A1 = CLBLL_L_X100Y133_SLICE_X156Y133_A5Q;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_A6 = CLBLM_L_X98Y130_SLICE_X154Y130_A5Q;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A3 = CLBLM_L_X98Y111_SLICE_X155Y111_C5Q;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A4 = CLBLM_L_X98Y111_SLICE_X155Y111_A5Q;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_A6 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_B6 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_C6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B3 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B4 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_B5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_C6 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_D6 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X156Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D1 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D3 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D4 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_D6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X155Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A2 = CLBLM_L_X98Y112_SLICE_X154Y112_A5Q;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A3 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A4 = CLBLL_L_X100Y111_SLICE_X156Y111_AQ;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_A6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_A6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B3 = CLBLM_L_X98Y112_SLICE_X155Y112_A5Q;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_B4 = CLBLM_R_X97Y112_SLICE_X152Y112_B5Q;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_B6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C1 = CLBLL_L_X100Y112_SLICE_X156Y112_CO6;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_C2 = CLBLL_L_X100Y112_SLICE_X157Y112_A5Q;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_C6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D1 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D2 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D3 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D4 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D5 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_D6 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D1 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D2 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D3 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D4 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D5 = 1'b1;
  assign CLBLL_L_X100Y130_SLICE_X157Y130_D6 = 1'b1;
  assign CLBLM_L_X98Y112_SLICE_X154Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A5 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A6 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_B1 = 1'b1;
  assign LIOI3_X0Y241_OLOGIC_X0Y241_D1 = 1'b0;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A2 = CLBLM_R_X101Y127_SLICE_X159Y127_A5Q;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A3 = CLBLM_R_X101Y126_SLICE_X159Y126_AQ;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A4 = CLBLM_L_X98Y125_SLICE_X155Y125_A5Q;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A5 = CLBLL_L_X100Y124_SLICE_X156Y124_AQ;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_A6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B1 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B2 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B3 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B4 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B5 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_B6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C1 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C2 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C3 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C4 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C5 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_C6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D1 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D2 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D3 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D4 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D5 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_D6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X159Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A2 = CLBLM_R_X101Y126_SLICE_X158Y126_A5Q;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A3 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A4 = CLBLM_R_X103Y125_SLICE_X162Y125_AQ;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A5 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_A6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B3 = CLBLL_L_X100Y124_SLICE_X157Y124_B5Q;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B4 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C1 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C2 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C3 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C4 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C5 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_C6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D1 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D2 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D3 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D4 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D5 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_D6 = 1'b1;
  assign CLBLM_R_X101Y126_SLICE_X158Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A1 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A2 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A3 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A4 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A5 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_A6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = 1'b0;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B1 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B2 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B3 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B4 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B5 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_B6 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C1 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C2 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C3 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C4 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C5 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_C6 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D1 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D2 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D3 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D4 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D5 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X155Y113_D6 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A2 = CLBLM_R_X97Y113_SLICE_X152Y113_A5Q;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A3 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A4 = CLBLM_L_X98Y113_SLICE_X154Y113_BO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A5 = CLBLM_L_X98Y112_SLICE_X154Y112_B5Q;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_A6 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B1 = CLBLL_L_X100Y113_SLICE_X156Y113_DO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B2 = CLBLL_L_X100Y113_SLICE_X156Y113_C5Q;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B5 = CLBLM_L_X98Y112_SLICE_X154Y112_AQ;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_B6 = CLBLM_R_X95Y116_SLICE_X150Y116_CO6;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B3 = CLBLL_L_X102Y127_SLICE_X160Y127_C5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C1 = CLBLM_L_X98Y115_SLICE_X154Y115_AQ;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C2 = CLBLL_L_X100Y113_SLICE_X157Y113_A5Q;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C4 = CLBLM_R_X95Y113_SLICE_X151Y113_DO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_C6 = CLBLM_L_X98Y114_SLICE_X154Y114_DO6;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D1 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D2 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D3 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D4 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D5 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_D6 = 1'b1;
  assign CLBLM_L_X98Y113_SLICE_X154Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_C1 = CLBLM_L_X90Y129_SLICE_X142Y129_AQ;
  assign RIOB33_X105Y183_IOB_X1Y184_O = 1'b0;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = 1'b0;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C4 = CLBLM_R_X95Y119_SLICE_X150Y119_BQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = 1'b0;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A2 = CLBLL_L_X100Y129_SLICE_X156Y129_AQ;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A3 = CLBLM_R_X101Y127_SLICE_X159Y127_AQ;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A4 = CLBLM_L_X98Y126_SLICE_X155Y126_A5Q;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A5 = CLBLM_R_X97Y126_SLICE_X153Y126_AQ;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_A6 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_D1 = CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B1 = CLBLL_L_X102Y127_SLICE_X160Y127_CQ;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B3 = CLBLM_R_X101Y127_SLICE_X159Y127_AQ;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B4 = CLBLL_L_X102Y129_SLICE_X160Y129_CQ;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B5 = CLBLL_L_X102Y127_SLICE_X160Y127_C5Q;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_B6 = CLBLL_L_X102Y127_SLICE_X160Y127_BQ;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_T1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C2 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C3 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_C6 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_D1 = CLBLL_L_X102Y117_SLICE_X160Y117_CO6;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B5 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D2 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D3 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D5 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_D6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A5 = CLBLM_R_X101Y136_SLICE_X158Y136_A5Q;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A6 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X159Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_T1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A2 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A3 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D3 = CLBLM_R_X95Y119_SLICE_X150Y119_BQ;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_A6 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B2 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B3 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B5 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_B6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_C1 = CLBLL_L_X100Y124_SLICE_X157Y124_CO6;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C2 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C3 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_C6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B2 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C5 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D1 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D2 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D3 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D4 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D5 = 1'b1;
  assign CLBLM_R_X101Y127_SLICE_X158Y127_D6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B6 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A1 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A2 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A3 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A4 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A5 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_A6 = 1'b1;
  assign CLBLL_L_X100Y125_SLICE_X157Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B1 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B2 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B3 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B4 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B5 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C1 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C1 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C2 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C3 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C4 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C5 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_C6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C2 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D1 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C3 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D2 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D1 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D2 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D3 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D4 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D5 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X155Y114_D6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C6 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A2 = CLBLM_L_X98Y113_SLICE_X154Y113_A5Q;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A3 = CLBLM_R_X95Y115_SLICE_X150Y115_A5Q;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A4 = CLBLL_L_X100Y114_SLICE_X156Y114_CO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A5 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_A6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_C5 = CLBLM_R_X89Y122_SLICE_X140Y122_DO6;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B2 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B3 = CLBLM_L_X98Y115_SLICE_X154Y115_B5Q;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B4 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B5 = CLBLM_R_X97Y115_SLICE_X153Y115_AQ;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_B6 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C1 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C2 = CLBLM_L_X98Y114_SLICE_X154Y114_CQ;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C4 = CLBLM_L_X98Y114_SLICE_X154Y114_BQ;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C5 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_C6 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D1 = CLBLM_L_X98Y114_SLICE_X154Y114_C5Q;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D2 = CLBLM_L_X98Y114_SLICE_X154Y114_CQ;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D3 = CLBLM_R_X97Y115_SLICE_X153Y115_AQ;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D4 = CLBLM_L_X98Y114_SLICE_X154Y114_BQ;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_D6 = 1'b1;
  assign CLBLM_L_X98Y114_SLICE_X154Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D3 = 1'b1;
  assign CLBLM_R_X93Y121_SLICE_X146Y121_D1 = CLBLM_L_X92Y121_SLICE_X144Y121_BQ;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D5 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A2 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A5 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_A6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B2 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B5 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_B6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C2 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C5 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_C6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D2 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D5 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X159Y128_D6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A2 = CLBLM_R_X101Y129_SLICE_X158Y129_B5Q;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A3 = CLBLL_L_X100Y129_SLICE_X157Y129_A5Q;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A5 = CLBLL_L_X100Y126_SLICE_X157Y126_DO6;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_A6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B2 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B5 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_B6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C2 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C3 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C4 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C5 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_C6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A2 = CLBLM_R_X97Y133_SLICE_X152Y133_A5Q;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A3 = CLBLL_L_X100Y133_SLICE_X156Y133_AQ;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A4 = CLBLM_L_X98Y132_SLICE_X154Y132_A5Q;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A5 = CLBLL_L_X100Y134_SLICE_X156Y134_B5Q;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_A6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D1 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B5 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_B6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_D6 = 1'b1;
  assign CLBLM_R_X101Y128_SLICE_X158Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C5 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_C6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A2 = CLBLM_R_X97Y115_SLICE_X152Y115_AQ;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A3 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A4 = CLBLM_L_X98Y115_SLICE_X155Y115_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A5 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_A6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B2 = CLBLM_L_X98Y115_SLICE_X155Y115_BQ;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D5 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_D6 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X156Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B3 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B4 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B5 = CLBLM_L_X98Y114_SLICE_X154Y114_AQ;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_B6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C1 = CLBLM_L_X98Y115_SLICE_X155Y115_C5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C2 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C4 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C5 = CLBLM_L_X90Y115_SLICE_X143Y115_AQ;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_C6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D2 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D3 = CLBLM_L_X98Y115_SLICE_X155Y115_BQ;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D4 = CLBLM_L_X98Y115_SLICE_X155Y115_A5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D5 = CLBLM_L_X98Y115_SLICE_X155Y115_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_D6 = CLBLM_L_X98Y114_SLICE_X154Y114_AQ;
  assign CLBLM_L_X98Y115_SLICE_X155Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A5 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_A6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A2 = CLBLM_L_X98Y115_SLICE_X155Y115_CQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A5 = CLBLM_L_X98Y115_SLICE_X154Y115_A5Q;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B5 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B2 = CLBLM_L_X98Y115_SLICE_X154Y115_BQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B3 = CLBLM_R_X97Y116_SLICE_X152Y116_AQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_B6 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C5 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_C6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C4 = CLBLM_L_X98Y115_SLICE_X154Y115_A5Q;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C5 = CLBLM_L_X98Y115_SLICE_X154Y115_DO6;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C6 = CLBLL_L_X100Y115_SLICE_X156Y115_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_C3 = CLBLM_R_X95Y115_SLICE_X150Y115_DO6;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D1 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D2 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D3 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D4 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D5 = 1'b1;
  assign CLBLL_L_X100Y133_SLICE_X157Y133_D6 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D2 = 1'b1;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D3 = CLBLM_R_X97Y116_SLICE_X152Y116_AQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D4 = CLBLM_L_X98Y115_SLICE_X154Y115_BQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D5 = CLBLM_L_X98Y115_SLICE_X154Y115_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_D6 = CLBLM_L_X98Y114_SLICE_X154Y114_B5Q;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_D1 = CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  assign LIOB33_X0Y59_IOB_X0Y60_T = 1'b1;
  assign LIOB33_X0Y59_IOB_X0Y59_T = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A1 = CLBLL_L_X102Y129_SLICE_X160Y129_A5Q;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A4 = CLBLM_R_X101Y129_SLICE_X159Y129_BO6;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A5 = CLBLM_R_X101Y129_SLICE_X158Y129_DO6;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_A6 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B3 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B4 = CLBLL_L_X100Y129_SLICE_X157Y129_A5Q;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B5 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C1 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C2 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C3 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C4 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C5 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_C6 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D1 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D2 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D3 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D4 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D5 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_D6 = 1'b1;
  assign LIOI3_X0Y241_OLOGIC_X0Y242_D1 = 1'b0;
  assign CLBLM_R_X101Y129_SLICE_X159Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A2 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A3 = CLBLM_R_X101Y129_SLICE_X158Y129_AQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A4 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A5 = CLBLM_R_X101Y129_SLICE_X159Y129_AQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_A6 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B2 = CLBLM_R_X101Y129_SLICE_X158Y129_BQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B3 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B4 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B5 = CLBLM_R_X101Y130_SLICE_X158Y130_CQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_B6 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C1 = CLBLM_R_X101Y129_SLICE_X158Y129_BQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C2 = CLBLM_R_X101Y130_SLICE_X158Y130_BQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C4 = CLBLM_R_X101Y130_SLICE_X158Y130_CQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C5 = CLBLM_R_X101Y129_SLICE_X158Y129_B5Q;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_C6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = 1'b0;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A1 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A2 = CLBLM_R_X101Y134_SLICE_X158Y134_AQ;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A3 = CLBLL_L_X100Y134_SLICE_X156Y134_AQ;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A5 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_A6 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D1 = CLBLM_R_X101Y129_SLICE_X159Y129_AQ;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B1 = CLBLM_R_X97Y133_SLICE_X153Y133_A5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B2 = CLBLL_L_X100Y134_SLICE_X156Y134_BQ;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B3 = CLBLM_L_X98Y134_SLICE_X154Y134_A5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B5 = CLBLM_L_X98Y132_SLICE_X155Y132_C5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_B6 = 1'b1;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D2 = CLBLM_R_X101Y129_SLICE_X158Y129_AQ;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y129_SLICE_X158Y129_D4 = CLBLM_R_X101Y129_SLICE_X158Y129_A5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C1 = CLBLM_L_X98Y132_SLICE_X155Y132_C5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C2 = CLBLM_R_X101Y134_SLICE_X158Y134_AQ;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C3 = CLBLL_L_X100Y134_SLICE_X156Y134_AQ;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C4 = CLBLL_L_X100Y134_SLICE_X156Y134_A5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_C6 = CLBLM_R_X101Y134_SLICE_X159Y134_BQ;
  assign CLBLM_L_X94Y118_SLICE_X149Y118_B4 = CLBLM_R_X93Y114_SLICE_X146Y114_B5Q;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A2 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A3 = CLBLM_L_X92Y116_SLICE_X145Y116_A5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A4 = CLBLM_R_X97Y116_SLICE_X153Y116_B5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A6 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D1 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D2 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D3 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D4 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D5 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_D6 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_A5 = CLBLL_L_X100Y116_SLICE_X156Y116_CO6;
  assign CLBLL_L_X100Y134_SLICE_X156Y134_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B2 = CLBLM_L_X98Y116_SLICE_X155Y116_BQ;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B3 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B4 = CLBLL_L_X100Y117_SLICE_X156Y117_A5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B5 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_B6 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C1 = CLBLM_L_X98Y115_SLICE_X155Y115_C5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C3 = CLBLM_L_X92Y116_SLICE_X144Y116_DO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C4 = CLBLM_L_X98Y116_SLICE_X155Y116_A5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C5 = CLBLM_L_X98Y116_SLICE_X155Y116_DO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_T1 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_D1 = CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D1 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D2 = CLBLM_R_X97Y116_SLICE_X153Y116_B5Q;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D4 = CLBLM_L_X98Y116_SLICE_X155Y116_BQ;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D5 = CLBLM_L_X98Y116_SLICE_X155Y116_B5Q;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A1 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A2 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A3 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A4 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A5 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_A6 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X155Y116_D6 = CLBLL_L_X100Y117_SLICE_X156Y117_A5Q;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A1 = CLBLL_L_X100Y116_SLICE_X157Y116_DO6;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A5 = CLBLL_L_X100Y114_SLICE_X156Y114_AQ;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_A6 = CLBLL_L_X100Y116_SLICE_X157Y116_B5Q;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B1 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B2 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B3 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B4 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B5 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_B6 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C1 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C2 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C3 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C4 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C5 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_C6 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B1 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B2 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B3 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B4 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B5 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_B6 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D1 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D2 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D3 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D4 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D5 = 1'b1;
  assign CLBLL_L_X100Y134_SLICE_X157Y134_D6 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C4 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C5 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D1 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D2 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D3 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D4 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D5 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = 1'b0;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C1 = 1'b1;
  assign LIOI3_X0Y241_OLOGIC_X0Y241_T1 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C2 = 1'b1;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C3 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A5 = CLBLM_L_X92Y119_SLICE_X145Y119_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y116_SLICE_X154Y116_C6 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y184_T = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y183_T = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B5 = CLBLM_L_X92Y120_SLICE_X145Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B6 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A3 = CLBLM_R_X101Y131_SLICE_X159Y131_DQ;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C2 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A5 = CLBLM_R_X101Y130_SLICE_X159Y130_CO6;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B2 = CLBLM_R_X101Y130_SLICE_X159Y130_BQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B3 = CLBLM_R_X101Y130_SLICE_X159Y130_AQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B4 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B5 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = 1'b0;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C1 = CLBLL_L_X102Y130_SLICE_X160Y130_AQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C2 = CLBLM_R_X101Y131_SLICE_X159Y131_A5Q;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C3 = CLBLM_R_X101Y130_SLICE_X159Y130_BQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C4 = CLBLM_R_X101Y130_SLICE_X159Y130_AQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C5 = CLBLM_R_X101Y130_SLICE_X159Y130_B5Q;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y132_SLICE_X153Y132_D6 = CLBLM_L_X98Y133_SLICE_X155Y133_BQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D1 = CLBLM_L_X98Y131_SLICE_X155Y131_DQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D3 = CLBLM_R_X101Y130_SLICE_X159Y130_BQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D4 = CLBLM_R_X101Y130_SLICE_X159Y130_AQ;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D5 = CLBLM_R_X101Y130_SLICE_X159Y130_B5Q;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_D6 = CLBLM_R_X101Y131_SLICE_X159Y131_A5Q;
  assign CLBLM_R_X101Y130_SLICE_X159Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A2 = CLBLM_R_X101Y130_SLICE_X158Y130_A5Q;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A3 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A4 = CLBLL_L_X102Y130_SLICE_X160Y130_AQ;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A5 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_A6 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B1 = CLBLM_R_X101Y130_SLICE_X158Y130_DO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B2 = CLBLM_R_X101Y129_SLICE_X158Y129_CO6;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B5 = CLBLL_L_X102Y129_SLICE_X160Y129_AQ;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_B6 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C1 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C2 = CLBLM_R_X101Y129_SLICE_X158Y129_A5Q;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C3 = CLBLM_R_X101Y130_SLICE_X158Y130_BQ;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C5 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D5 = 1'b1;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_D6 = CLBLM_R_X101Y128_SLICE_X158Y128_A5Q;
  assign CLBLM_R_X101Y130_SLICE_X158Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A2 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A3 = CLBLM_L_X98Y117_SLICE_X155Y117_AQ;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A4 = CLBLL_L_X100Y114_SLICE_X156Y114_AQ;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A5 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_A6 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B2 = CLBLM_L_X98Y117_SLICE_X155Y117_BQ;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B3 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B4 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B5 = CLBLM_L_X94Y116_SLICE_X149Y116_AQ;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_B6 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C1 = CLBLM_L_X98Y117_SLICE_X155Y117_DO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C2 = CLBLL_L_X100Y118_SLICE_X157Y118_A5Q;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C3 = CLBLM_R_X93Y117_SLICE_X146Y117_CO6;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_C6 = CLBLM_L_X98Y117_SLICE_X155Y117_AQ;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_C5 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D1 = CLBLM_L_X94Y116_SLICE_X149Y116_AQ;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D3 = CLBLM_L_X98Y119_SLICE_X155Y119_B5Q;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D4 = CLBLM_L_X98Y117_SLICE_X155Y117_BQ;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D5 = CLBLM_L_X98Y117_SLICE_X155Y117_B5Q;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_D6 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X155Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A1 = CLBLM_R_X97Y117_SLICE_X153Y117_BQ;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A2 = CLBLM_R_X97Y118_SLICE_X153Y118_BQ;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A4 = CLBLM_R_X97Y117_SLICE_X153Y117_C5Q;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A5 = CLBLL_L_X100Y118_SLICE_X157Y118_C5Q;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_A6 = CLBLM_R_X97Y117_SLICE_X152Y117_B5Q;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B1 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B2 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B3 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B4 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B5 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_B6 = 1'b1;
  assign CLBLM_L_X90Y122_SLICE_X143Y122_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C1 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C2 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C3 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C4 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C5 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_C6 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D1 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D2 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D3 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D4 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D5 = 1'b1;
  assign CLBLM_L_X98Y117_SLICE_X154Y117_D6 = 1'b1;
  assign CLBLL_L_X100Y120_SLICE_X156Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C2 = CLBLM_L_X90Y120_SLICE_X143Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C3 = CLBLM_R_X93Y124_SLICE_X147Y124_DO6;
  assign CLBLM_L_X90Y120_SLICE_X143Y120_D3 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C5 = CLBLM_L_X92Y120_SLICE_X144Y120_DO6;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A1 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A2 = CLBLM_R_X101Y130_SLICE_X159Y130_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A3 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A5 = CLBLM_R_X101Y131_SLICE_X158Y131_AQ;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_A6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B1 = CLBLM_R_X101Y132_SLICE_X159Y132_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B2 = CLBLL_L_X102Y131_SLICE_X160Y131_AQ;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B3 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B5 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_B6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C1 = CLBLM_R_X101Y133_SLICE_X159Y133_AQ;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C3 = CLBLM_R_X101Y128_SLICE_X158Y128_A5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C4 = CLBLL_L_X102Y131_SLICE_X160Y131_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C5 = CLBLM_R_X101Y131_SLICE_X159Y131_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_C6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D1 = CLBLM_R_X101Y131_SLICE_X159Y131_DQ;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D3 = CLBLM_R_X101Y131_SLICE_X158Y131_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D4 = CLBLM_R_X101Y131_SLICE_X159Y131_A5Q;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D5 = CLBLM_R_X101Y131_SLICE_X159Y131_CQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A2 = CLBLM_R_X95Y113_SLICE_X150Y113_BQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A3 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A4 = CLBLM_R_X95Y113_SLICE_X151Y113_B5Q;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A5 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_A6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X159Y131_D6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B2 = CLBLM_R_X95Y111_SLICE_X151Y111_BQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B3 = CLBLM_R_X95Y111_SLICE_X151Y111_AQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B4 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B5 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_B6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A2 = CLBLM_R_X101Y131_SLICE_X159Y131_D5Q;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A3 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C1 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C2 = CLBLM_R_X95Y113_SLICE_X150Y113_BQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C3 = CLBLM_R_X95Y111_SLICE_X151Y111_BQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C5 = CLBLM_R_X95Y111_SLICE_X151Y111_B5Q;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_C6 = CLBLM_R_X95Y111_SLICE_X151Y111_AQ;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B2 = CLBLM_R_X101Y131_SLICE_X158Y131_BQ;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_B3 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C2 = CLBLM_R_X101Y131_SLICE_X158Y131_AQ;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C3 = CLBLM_R_X101Y130_SLICE_X158Y130_A5Q;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C4 = CLBLM_R_X101Y131_SLICE_X158Y131_BQ;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D1 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D2 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D3 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D4 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D5 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_D6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C5 = CLBLM_R_X101Y131_SLICE_X158Y131_B5Q;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y111_SLICE_X151Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D1 = CLBLM_R_X101Y131_SLICE_X159Y131_AQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A1 = CLBLM_R_X95Y112_SLICE_X150Y112_DO6;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A2 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A3 = CLBLM_R_X97Y111_SLICE_X152Y111_A5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A5 = CLBLM_R_X95Y111_SLICE_X150Y111_C5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_A6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D2 = CLBLM_R_X101Y131_SLICE_X158Y131_AQ;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D3 = CLBLM_L_X98Y131_SLICE_X155Y131_D5Q;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D4 = CLBLM_R_X101Y131_SLICE_X158Y131_BQ;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_D5 = CLBLM_R_X101Y131_SLICE_X158Y131_B5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B1 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B3 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B4 = CLBLM_L_X94Y111_SLICE_X149Y111_B5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B5 = CLBLM_L_X94Y112_SLICE_X149Y112_BQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_B6 = 1'b1;
  assign CLBLM_R_X101Y131_SLICE_X158Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C1 = CLBLM_R_X95Y111_SLICE_X150Y111_BQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C2 = CLBLM_R_X95Y111_SLICE_X150Y111_CQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C3 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C5 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_C6 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D1 = CLBLM_R_X95Y111_SLICE_X150Y111_BQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D2 = CLBLM_R_X95Y111_SLICE_X150Y111_CQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D3 = CLBLM_R_X95Y111_SLICE_X150Y111_C5Q;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D4 = 1'b1;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D5 = CLBLM_L_X94Y112_SLICE_X149Y112_BQ;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y111_SLICE_X150Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y51_IOB_X0Y52_O = 1'b0;
  assign LIOB33_X0Y51_IOB_X0Y51_O = 1'b0;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = 1'b0;
  assign LIOB33_X0Y51_IOB_X0Y52_T = 1'b1;
  assign LIOB33_X0Y51_IOB_X0Y51_T = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = 1'b0;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_D1 = CLBLL_L_X102Y116_SLICE_X160Y116_AO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_T1 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_D1 = CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_T1 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = 1'b0;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C4 = CLBLM_R_X95Y120_SLICE_X150Y120_BQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = 1'b0;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C5 = CLBLM_R_X95Y120_SLICE_X150Y120_B5Q;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C6 = CLBLM_R_X95Y122_SLICE_X150Y122_BQ;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A3 = CLBLM_R_X101Y131_SLICE_X159Y131_C5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A4 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A5 = CLBLM_R_X101Y132_SLICE_X159Y132_CO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B3 = CLBLM_R_X101Y132_SLICE_X159Y132_AQ;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B4 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B5 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_B2 = CLBLM_R_X101Y132_SLICE_X159Y132_BQ;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B4 = CLBLL_L_X100Y126_SLICE_X156Y126_DO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C2 = CLBLM_R_X101Y131_SLICE_X159Y131_B5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C3 = CLBLM_R_X101Y132_SLICE_X159Y132_BQ;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C4 = CLBLM_R_X101Y132_SLICE_X159Y132_AQ;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C5 = CLBLM_R_X101Y132_SLICE_X159Y132_B5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_C6 = CLBLM_R_X101Y132_SLICE_X158Y132_A5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D1 = CLBLM_L_X98Y130_SLICE_X155Y130_D5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D2 = CLBLM_R_X101Y131_SLICE_X159Y131_B5Q;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D3 = CLBLM_R_X101Y132_SLICE_X159Y132_BQ;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D4 = CLBLM_R_X101Y132_SLICE_X159Y132_AQ;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D5 = CLBLM_R_X101Y132_SLICE_X159Y132_B5Q;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A1 = CLBLM_R_X93Y114_SLICE_X147Y114_CO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A4 = CLBLM_R_X97Y112_SLICE_X152Y112_A5Q;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A5 = CLBLM_R_X95Y113_SLICE_X151Y113_AQ;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B6 = CLBLM_L_X92Y127_SLICE_X145Y127_CO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_A6 = CLBLM_R_X95Y111_SLICE_X151Y111_CO6;
  assign CLBLM_R_X101Y132_SLICE_X159Y132_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B1 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B2 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B3 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B4 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B5 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_B6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A2 = CLBLM_R_X101Y132_SLICE_X158Y132_A5Q;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A3 = CLBLM_R_X101Y130_SLICE_X158Y130_AQ;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_A4 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C1 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C2 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C3 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C4 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C5 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_C6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B1 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B2 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B3 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C1 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B4 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_B5 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C5 = CLBLL_L_X100Y124_SLICE_X157Y124_DO6;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D1 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D2 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D3 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D4 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_C6 = CLBLM_R_X101Y126_SLICE_X158Y126_AQ;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D5 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X151Y112_D6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_C6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D1 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A1 = CLBLM_R_X95Y113_SLICE_X150Y113_CO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A3 = CLBLM_R_X95Y112_SLICE_X150Y112_B5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A4 = CLBLM_R_X93Y111_SLICE_X147Y111_B5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A5 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_A6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D2 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D3 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D4 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_D5 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B2 = CLBLM_R_X93Y111_SLICE_X147Y111_A5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B3 = CLBLM_R_X95Y111_SLICE_X150Y111_A5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B4 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B5 = CLBLM_R_X95Y112_SLICE_X150Y112_CO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_B6 = 1'b1;
  assign CLBLM_R_X101Y132_SLICE_X158Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A3 = CLBLM_L_X98Y119_SLICE_X154Y119_A5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A4 = CLBLL_L_X100Y119_SLICE_X156Y119_AO6;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A5 = CLBLM_L_X92Y118_SLICE_X144Y118_BO6;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C2 = CLBLM_R_X95Y113_SLICE_X150Y113_A5Q;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B2 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B3 = CLBLM_L_X98Y119_SLICE_X155Y119_AQ;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B4 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B5 = CLBLM_L_X98Y117_SLICE_X155Y117_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_B6 = 1'b1;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C1 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C2 = CLBLM_L_X98Y119_SLICE_X155Y119_CQ;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C4 = CLBLM_R_X97Y119_SLICE_X152Y119_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C5 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_C6 = 1'b1;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D4 = CLBLM_R_X93Y112_SLICE_X146Y112_CO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_D3 = CLBLL_L_X102Y126_SLICE_X160Y126_DO6;
  assign CLBLM_R_X95Y112_SLICE_X150Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D1 = CLBLM_L_X98Y119_SLICE_X155Y119_C5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D2 = CLBLM_L_X98Y119_SLICE_X155Y119_CQ;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D3 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D4 = CLBLM_L_X98Y120_SLICE_X155Y120_A5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D5 = CLBLM_R_X97Y119_SLICE_X152Y119_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_C1 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D1 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X155Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y53_IOB_X0Y53_O = 1'b0;
  assign LIOB33_X0Y53_IOB_X0Y54_T = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A2 = CLBLM_L_X98Y119_SLICE_X154Y119_A5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A3 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A4 = CLBLM_R_X97Y122_SLICE_X152Y122_AQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A5 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_A6 = 1'b1;
  assign LIOB33_X0Y53_IOB_X0Y53_T = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B2 = CLBLM_L_X90Y118_SLICE_X142Y118_CO6;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B3 = CLBLM_L_X98Y119_SLICE_X154Y119_AQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_B6 = CLBLM_L_X98Y119_SLICE_X154Y119_CO6;
  assign CLBLL_L_X100Y126_SLICE_X157Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_BX = CLBLM_L_X98Y119_SLICE_X154Y119_CO5;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C1 = CLBLM_L_X98Y120_SLICE_X154Y120_CQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C2 = CLBLM_L_X98Y119_SLICE_X154Y119_B5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C3 = CLBLM_R_X97Y118_SLICE_X153Y118_C5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C5 = CLBLM_L_X98Y119_SLICE_X154Y119_BQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_C6 = 1'b1;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y122_SLICE_X146Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D1 = CLBLM_L_X98Y120_SLICE_X154Y120_CQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D3 = CLBLM_R_X97Y118_SLICE_X153Y118_C5Q;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D4 = CLBLL_L_X100Y118_SLICE_X157Y118_BQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D5 = CLBLM_L_X98Y119_SLICE_X154Y119_BQ;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_D6 = CLBLM_L_X98Y119_SLICE_X154Y119_B5Q;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1 = 1'b0;
  assign CLBLM_L_X98Y119_SLICE_X154Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y117_IOB_X0Y118_T = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_T = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_T1 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A1 = CLBLL_L_X100Y134_SLICE_X156Y134_A5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A2 = CLBLM_R_X101Y134_SLICE_X158Y134_A5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A4 = CLBLM_R_X101Y131_SLICE_X159Y131_D5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A5 = CLBLM_R_X101Y131_SLICE_X159Y131_C5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_A6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B1 = CLBLM_R_X101Y135_SLICE_X159Y135_A5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B2 = CLBLM_R_X101Y134_SLICE_X159Y134_CQ;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B4 = CLBLL_L_X100Y133_SLICE_X156Y133_AQ;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B5 = CLBLM_R_X101Y134_SLICE_X159Y134_AQ;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_B6 = CLBLM_R_X101Y134_SLICE_X159Y134_C5Q;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C1 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C2 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C3 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C4 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C5 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_C6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D1 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D2 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D3 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D4 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D5 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A1 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A2 = CLBLM_R_X95Y113_SLICE_X151Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A4 = CLBLM_R_X95Y116_SLICE_X151Y116_AQ;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A5 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_A6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X159Y133_D6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B1 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B2 = CLBLM_R_X95Y113_SLICE_X151Y113_BQ;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B4 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B5 = CLBLM_R_X95Y114_SLICE_X150Y114_AQ;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_B6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C3 = CLBLM_L_X94Y113_SLICE_X149Y113_CO6;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C4 = CLBLM_R_X95Y113_SLICE_X151Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C5 = CLBLM_R_X95Y113_SLICE_X151Y113_DO6;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_C6 = CLBLM_R_X97Y112_SLICE_X153Y112_B5Q;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B2 = CLBLM_R_X101Y133_SLICE_X158Y133_BQ;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B3 = CLBLM_R_X101Y133_SLICE_X158Y133_AQ;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B4 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_B5 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D1 = CLBLM_R_X95Y114_SLICE_X150Y114_AQ;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D2 = CLBLM_R_X95Y111_SLICE_X151Y111_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D3 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D4 = CLBLM_R_X95Y113_SLICE_X151Y113_BQ;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D5 = CLBLM_R_X95Y113_SLICE_X151Y113_B5Q;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C3 = CLBLM_R_X101Y133_SLICE_X158Y133_BQ;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y113_SLICE_X151Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D1 = CLBLM_L_X98Y132_SLICE_X155Y132_CQ;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D2 = CLBLM_R_X101Y133_SLICE_X158Y133_AQ;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A1 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A2 = CLBLM_R_X95Y113_SLICE_X150Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A3 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A4 = CLBLM_R_X97Y111_SLICE_X153Y111_AQ;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_A6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D3 = CLBLM_R_X101Y134_SLICE_X158Y134_A5Q;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D4 = CLBLM_R_X101Y133_SLICE_X158Y133_BQ;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D5 = CLBLM_R_X101Y133_SLICE_X158Y133_B5Q;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B1 = CLBLM_R_X95Y114_SLICE_X150Y114_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B2 = CLBLM_L_X94Y113_SLICE_X149Y113_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B3 = CLBLM_R_X95Y112_SLICE_X151Y112_AO6;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B4 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_B6 = 1'b1;
  assign CLBLM_R_X101Y133_SLICE_X158Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A2 = CLBLM_R_X101Y118_SLICE_X158Y118_A5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A3 = CLBLM_L_X98Y119_SLICE_X155Y119_C5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A4 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A5 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_A6 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D6 = CLBLM_R_X89Y124_SLICE_X141Y124_BQ;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_C2 = CLBLM_R_X95Y113_SLICE_X150Y113_AQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B2 = CLBLM_L_X98Y120_SLICE_X155Y120_BQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B3 = CLBLM_L_X98Y120_SLICE_X155Y120_AQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B4 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B5 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_B6 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D1 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C1 = CLBLM_L_X98Y120_SLICE_X154Y120_AQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C2 = CLBLM_L_X98Y121_SLICE_X154Y121_DQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C4 = CLBLM_R_X101Y119_SLICE_X158Y119_CQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C5 = CLBLM_L_X98Y120_SLICE_X154Y120_C5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_C6 = CLBLM_L_X98Y120_SLICE_X154Y120_A5Q;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D2 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D3 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D4 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D5 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_D6 = 1'b1;
  assign CLBLM_R_X95Y113_SLICE_X150Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D1 = CLBLM_L_X98Y120_SLICE_X155Y120_BQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D2 = CLBLM_L_X98Y120_SLICE_X155Y120_AQ;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D4 = CLBLM_R_X101Y118_SLICE_X158Y118_A5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D5 = CLBLM_L_X98Y120_SLICE_X155Y120_B5Q;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_D6 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X155Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A2 = CLBLM_R_X97Y122_SLICE_X152Y122_AQ;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A4 = CLBLM_L_X98Y120_SLICE_X154Y120_BO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A5 = CLBLM_R_X89Y120_SLICE_X140Y120_DO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_AX = CLBLM_L_X98Y120_SLICE_X154Y120_BO5;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B2 = CLBLM_L_X98Y120_SLICE_X154Y120_A5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B3 = CLBLM_L_X98Y120_SLICE_X154Y120_AQ;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B4 = CLBLM_L_X98Y121_SLICE_X154Y121_DQ;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B5 = CLBLM_L_X98Y120_SLICE_X154Y120_C5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_B6 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C1 = CLBLM_L_X98Y119_SLICE_X154Y119_BQ;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C2 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C4 = CLBLM_L_X98Y121_SLICE_X154Y121_DQ;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C5 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_C6 = 1'b1;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D3 = CLBLM_R_X103Y125_SLICE_X163Y125_DO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D4 = CLBLM_R_X97Y120_SLICE_X153Y120_B5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D5 = CLBLL_L_X100Y122_SLICE_X157Y122_B5Q;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_D6 = CLBLM_L_X98Y119_SLICE_X155Y119_DO6;
  assign CLBLM_L_X98Y120_SLICE_X154Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = 1'b0;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A1 = CLBLM_R_X101Y134_SLICE_X159Y134_DO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A3 = CLBLM_R_X101Y135_SLICE_X159Y135_DQ;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = 1'b0;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B2 = CLBLM_R_X101Y134_SLICE_X158Y134_BO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B3 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B5 = CLBLM_R_X101Y133_SLICE_X159Y133_A5Q;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C1 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C3 = CLBLM_R_X101Y134_SLICE_X159Y134_CQ;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C4 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C5 = CLBLM_R_X101Y134_SLICE_X159Y134_AQ;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_C6 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_D1 = CLBLL_L_X102Y119_SLICE_X160Y119_CO6;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D1 = CLBLM_R_X101Y134_SLICE_X159Y134_C5Q;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D2 = CLBLM_R_X101Y134_SLICE_X159Y134_CQ;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D3 = CLBLM_R_X101Y135_SLICE_X159Y135_A5Q;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D4 = CLBLM_R_X101Y134_SLICE_X159Y134_AQ;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A1 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A2 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A3 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A4 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A5 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_A6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X159Y134_D6 = CLBLL_L_X102Y134_SLICE_X160Y134_A5Q;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A1 = CLBLM_R_X101Y133_SLICE_X158Y133_B5Q;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B1 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B2 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B3 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B4 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B5 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A3 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_A4 = CLBLM_R_X101Y134_SLICE_X159Y134_BQ;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C1 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C2 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C3 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C4 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C5 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_C6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B1 = CLBLL_L_X100Y134_SLICE_X156Y134_A5Q;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B3 = CLBLM_R_X101Y134_SLICE_X158Y134_AQ;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B4 = CLBLM_R_X101Y134_SLICE_X159Y134_BQ;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B5 = CLBLM_R_X101Y132_SLICE_X158Y132_AQ;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_B6 = CLBLL_L_X100Y134_SLICE_X156Y134_AQ;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D1 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D2 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D3 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D4 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D5 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X151Y114_D6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C3 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C4 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_C6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D1 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A2 = CLBLM_R_X95Y114_SLICE_X150Y114_B5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A3 = CLBLM_R_X95Y113_SLICE_X151Y113_CO6;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A4 = CLBLM_R_X93Y120_SLICE_X147Y120_C5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A5 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_A6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D2 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D3 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D4 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_D5 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B2 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B3 = CLBLM_L_X94Y114_SLICE_X149Y114_BQ;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B4 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B5 = CLBLM_R_X95Y114_SLICE_X150Y114_C5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y134_SLICE_X158Y134_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A2 = CLBLM_L_X98Y121_SLICE_X155Y121_B5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A3 = CLBLM_L_X98Y121_SLICE_X155Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A4 = CLBLM_L_X98Y121_SLICE_X155Y121_AQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A5 = CLBLM_L_X98Y121_SLICE_X154Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_A6 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C1 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C2 = CLBLM_R_X95Y114_SLICE_X150Y114_CQ;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B2 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B3 = CLBLM_L_X98Y121_SLICE_X155Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B4 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B5 = CLBLM_L_X98Y123_SLICE_X155Y123_AQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_B6 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D1 = CLBLM_R_X95Y114_SLICE_X150Y114_C5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C1 = CLBLM_L_X98Y121_SLICE_X154Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C2 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C4 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C5 = CLBLL_L_X100Y121_SLICE_X157Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_C6 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D2 = CLBLM_R_X95Y114_SLICE_X150Y114_CQ;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D3 = CLBLM_R_X95Y115_SLICE_X150Y115_B5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D5 = CLBLM_R_X95Y114_SLICE_X150Y114_B5Q;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_D6 = 1'b1;
  assign CLBLM_R_X95Y114_SLICE_X150Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D1 = CLBLL_L_X102Y120_SLICE_X160Y120_D5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D2 = CLBLM_L_X98Y121_SLICE_X155Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D4 = CLBLM_L_X98Y121_SLICE_X154Y121_CQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D5 = CLBLM_L_X98Y121_SLICE_X155Y121_B5Q;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_D6 = CLBLM_L_X98Y121_SLICE_X155Y121_AQ;
  assign CLBLM_L_X98Y121_SLICE_X155Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A2 = CLBLM_L_X98Y121_SLICE_X154Y121_A5Q;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A3 = CLBLL_L_X100Y121_SLICE_X156Y121_AQ;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A4 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A5 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_A6 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B2 = CLBLM_L_X98Y121_SLICE_X154Y121_BQ;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B3 = CLBLM_L_X98Y121_SLICE_X154Y121_D5Q;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B4 = CLBLM_L_X98Y122_SLICE_X154Y122_BQ;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B5 = CLBLM_R_X97Y122_SLICE_X152Y122_BQ;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_B6 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C1 = CLBLM_L_X98Y121_SLICE_X154Y121_A5Q;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C5 = CLBLM_R_X93Y122_SLICE_X147Y122_DO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_C6 = CLBLM_L_X98Y121_SLICE_X155Y121_AO6;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D1 = CLBLM_L_X98Y120_SLICE_X154Y120_AQ;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D2 = CLBLM_L_X98Y122_SLICE_X154Y122_BQ;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D4 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D5 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_D6 = 1'b1;
  assign CLBLM_L_X98Y121_SLICE_X154Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A1 = CLBLM_L_X92Y121_SLICE_X145Y121_B5Q;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A2 = CLBLM_L_X92Y121_SLICE_X145Y121_BQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B1 = CLBLM_L_X92Y121_SLICE_X145Y121_BQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B3 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B4 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B5 = CLBLM_L_X92Y121_SLICE_X144Y121_CQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_B6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A2 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A3 = CLBLM_R_X101Y134_SLICE_X159Y134_C5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A4 = CLBLL_L_X102Y135_SLICE_X160Y135_AQ;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A5 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_A6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B2 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B3 = CLBLM_R_X101Y136_SLICE_X159Y136_B5Q;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C2 = CLBLM_L_X92Y121_SLICE_X145Y121_CQ;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B4 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B5 = CLBLL_L_X102Y136_SLICE_X160Y136_AQ;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_B6 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C3 = CLBLM_R_X93Y121_SLICE_X147Y121_AQ;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C1 = CLBLM_R_X101Y133_SLICE_X159Y133_A5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C2 = CLBLM_R_X101Y135_SLICE_X159Y135_CQ;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C3 = CLBLL_L_X102Y136_SLICE_X160Y136_B5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C5 = CLBLM_R_X101Y135_SLICE_X159Y135_B5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_C6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D1 = CLBLM_R_X101Y135_SLICE_X159Y135_C5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D2 = CLBLM_R_X101Y135_SLICE_X158Y135_A5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D3 = CLBLM_R_X101Y135_SLICE_X159Y135_DQ;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D5 = CLBLM_R_X101Y135_SLICE_X159Y135_A5Q;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A1 = CLBLM_R_X95Y114_SLICE_X150Y114_DO6;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A2 = CLBLM_R_X95Y115_SLICE_X150Y115_DO6;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A5 = CLBLM_R_X95Y116_SLICE_X151Y116_AQ;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_A6 = CLBLM_R_X97Y115_SLICE_X153Y115_A5Q;
  assign CLBLM_R_X101Y135_SLICE_X159Y135_D6 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B1 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B2 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B3 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B5 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_B6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A2 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_A3 = CLBLM_R_X101Y135_SLICE_X158Y135_AQ;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C1 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C2 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C3 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C5 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_C6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B2 = CLBLL_L_X102Y135_SLICE_X160Y135_AQ;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B3 = CLBLM_R_X101Y135_SLICE_X158Y135_AQ;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B4 = CLBLL_L_X100Y133_SLICE_X156Y133_A5Q;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B5 = CLBLM_R_X101Y135_SLICE_X159Y135_AQ;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_B6 = CLBLM_R_X101Y135_SLICE_X158Y135_A5Q;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D1 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D2 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D3 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D5 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X151Y115_D6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C3 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_A1 = CLBLM_L_X90Y122_SLICE_X142Y122_AQ;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_C6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D1 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A2 = CLBLM_R_X95Y116_SLICE_X150Y116_A5Q;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A3 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A5 = CLBLM_R_X93Y115_SLICE_X147Y115_AQ;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_A6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B2 = CLBLM_R_X95Y116_SLICE_X150Y116_BO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B3 = CLBLM_R_X95Y115_SLICE_X151Y115_AO6;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B4 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B5 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_B6 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A2 = CLBLM_L_X98Y122_SLICE_X155Y122_A5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A3 = CLBLM_R_X97Y124_SLICE_X152Y124_AQ;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A4 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A5 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_A6 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C1 = CLBLM_R_X97Y116_SLICE_X152Y116_BQ;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C2 = CLBLM_R_X95Y115_SLICE_X150Y115_CQ;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_C3 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B2 = CLBLM_L_X98Y122_SLICE_X155Y122_BQ;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B3 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B4 = CLBLL_L_X100Y123_SLICE_X156Y123_BQ;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B5 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_B6 = 1'b1;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D1 = CLBLM_R_X95Y115_SLICE_X150Y115_C5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C1 = CLBLM_L_X98Y122_SLICE_X155Y122_A5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C2 = CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C4 = CLBLM_R_X97Y122_SLICE_X152Y122_D5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C5 = CLBLM_L_X98Y122_SLICE_X155Y122_DO6;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D2 = CLBLM_R_X95Y115_SLICE_X150Y115_CQ;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D3 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D4 = CLBLM_R_X95Y115_SLICE_X150Y115_BQ;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D5 = CLBLM_R_X97Y116_SLICE_X152Y116_BQ;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y115_SLICE_X150Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D1 = CLBLM_L_X98Y122_SLICE_X155Y122_BQ;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D2 = CLBLM_R_X97Y122_SLICE_X153Y122_B5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D3 = CLBLL_L_X100Y123_SLICE_X156Y123_BQ;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D4 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D5 = CLBLM_L_X98Y122_SLICE_X155Y122_B5Q;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y122_SLICE_X155Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B5 = CLBLM_L_X90Y123_SLICE_X143Y123_C5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A2 = CLBLM_L_X98Y122_SLICE_X154Y122_A5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A3 = CLBLM_L_X98Y121_SLICE_X154Y121_AQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A4 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A5 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_A6 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_B6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C6 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B2 = CLBLM_L_X98Y123_SLICE_X154Y123_CQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B3 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B4 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B5 = CLBLM_R_X97Y122_SLICE_X152Y122_BQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_B6 = 1'b1;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C1 = CLBLM_R_X97Y122_SLICE_X152Y122_BQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C3 = CLBLM_L_X98Y122_SLICE_X154Y122_BQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C4 = CLBLM_L_X98Y121_SLICE_X154Y121_D5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C5 = CLBLM_R_X101Y123_SLICE_X159Y123_C5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_C6 = CLBLM_L_X98Y121_SLICE_X154Y121_BQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y123_SLICE_X143Y123_C2 = CLBLM_L_X90Y123_SLICE_X143Y123_CQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D2 = CLBLM_R_X97Y122_SLICE_X153Y122_AQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D3 = CLBLM_R_X101Y123_SLICE_X159Y123_CQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D4 = CLBLM_L_X98Y123_SLICE_X154Y123_CQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D5 = CLBLM_L_X98Y122_SLICE_X154Y122_B5Q;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_D6 = CLBLM_R_X97Y122_SLICE_X152Y122_CQ;
  assign CLBLM_L_X98Y122_SLICE_X154Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B1 = CLBLM_L_X92Y122_SLICE_X144Y122_DO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D1 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D2 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D3 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A5 = CLBLM_R_X101Y135_SLICE_X159Y135_CQ;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_A6 = CLBLM_R_X101Y136_SLICE_X159Y136_CO6;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B1 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B2 = CLBLM_R_X101Y136_SLICE_X159Y136_BQ;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B3 = CLBLM_R_X101Y136_SLICE_X159Y136_AQ;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B5 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_B6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C2 = CLBLM_R_X101Y136_SLICE_X158Y136_A5Q;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C3 = CLBLM_R_X101Y135_SLICE_X159Y135_B5Q;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C4 = CLBLM_R_X101Y136_SLICE_X159Y136_BQ;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C5 = CLBLM_R_X101Y136_SLICE_X159Y136_B5Q;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_C6 = CLBLM_R_X101Y136_SLICE_X159Y136_AQ;
  assign LIOB33_X0Y61_IOB_X0Y61_O = 1'b0;
  assign LIOB33_X0Y61_IOB_X0Y62_O = 1'b0;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y61_IOB_X0Y62_T = 1'b1;
  assign LIOB33_X0Y61_IOB_X0Y61_T = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D1 = CLBLL_L_X100Y134_SLICE_X156Y134_BQ;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D3 = CLBLM_R_X101Y135_SLICE_X159Y135_B5Q;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D4 = CLBLM_R_X101Y136_SLICE_X159Y136_BQ;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D5 = CLBLM_R_X101Y136_SLICE_X159Y136_B5Q;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A1 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A2 = CLBLM_R_X95Y116_SLICE_X151Y116_A5Q;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A4 = CLBLM_L_X90Y116_SLICE_X143Y116_AQ;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A5 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_A6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X159Y136_D6 = CLBLM_R_X101Y136_SLICE_X159Y136_AQ;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A1 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B1 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B2 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B3 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B4 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B5 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_B6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A3 = CLBLM_R_X101Y132_SLICE_X158Y132_AQ;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_A4 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C1 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C2 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C3 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C4 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B1 = CLBLM_L_X90Y123_SLICE_X142Y123_CQ;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C5 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_C6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B1 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_B2 = CLBLM_L_X90Y115_SLICE_X142Y115_A5Q;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B3 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B4 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_B5 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D1 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D2 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D3 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D4 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D5 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_D6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_C4 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A2 = CLBLL_L_X102Y128_SLICE_X161Y128_B5Q;
  assign CLBLM_R_X95Y116_SLICE_X151Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A1 = CLBLM_R_X95Y116_SLICE_X150Y116_AQ;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A3 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A2 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A3 = CLBLM_L_X94Y113_SLICE_X148Y113_AQ;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A4 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_A6 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D1 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D2 = 1'b1;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_D4 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B1 = CLBLM_R_X95Y114_SLICE_X150Y114_DO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B4 = CLBLM_R_X95Y114_SLICE_X150Y114_A5Q;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B5 = CLBLM_R_X95Y121_SLICE_X151Y121_CO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_B6 = CLBLM_L_X94Y116_SLICE_X149Y116_B5Q;
  assign CLBLM_R_X101Y136_SLICE_X158Y136_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = 1'b0;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A4 = CLBLM_L_X98Y123_SLICE_X155Y123_BO6;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A5 = CLBLM_L_X98Y121_SLICE_X154Y121_AQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_A6 = CLBLM_R_X93Y123_SLICE_X147Y123_DO6;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C1 = CLBLM_L_X94Y113_SLICE_X148Y113_AQ;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_AX = CLBLM_L_X98Y123_SLICE_X155Y123_BO5;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_C3 = CLBLM_R_X95Y116_SLICE_X150Y116_AQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B2 = CLBLM_L_X98Y123_SLICE_X155Y123_A5Q;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B3 = CLBLM_L_X98Y123_SLICE_X155Y123_AQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B4 = CLBLM_L_X98Y121_SLICE_X155Y121_BQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B5 = CLBLM_L_X98Y123_SLICE_X155Y123_C5Q;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_B6 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C1 = CLBLM_L_X98Y121_SLICE_X155Y121_BQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C2 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B1 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C4 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B2 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C5 = CLBLM_L_X98Y123_SLICE_X154Y123_AQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_C6 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D4 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B3 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_D6 = 1'b1;
  assign CLBLM_R_X95Y116_SLICE_X150Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D1 = CLBLM_L_X98Y123_SLICE_X155Y123_C5Q;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B4 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D4 = CLBLM_L_X98Y123_SLICE_X155Y123_A5Q;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D3 = CLBLL_L_X102Y124_SLICE_X160Y124_DQ;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B5 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D5 = CLBLM_L_X98Y123_SLICE_X155Y123_AQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_D6 = CLBLM_L_X98Y121_SLICE_X155Y121_BQ;
  assign CLBLM_L_X98Y123_SLICE_X155Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_D1 = 1'b0;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A4 = CLBLM_L_X98Y123_SLICE_X154Y123_BO6;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A5 = CLBLM_L_X98Y122_SLICE_X154Y122_A5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_A6 = CLBLM_R_X93Y123_SLICE_X146Y123_DO6;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_D1 = 1'b0;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_T1 = 1'b1;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_AX = CLBLM_L_X98Y123_SLICE_X154Y123_BO5;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_T1 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B2 = CLBLM_L_X98Y123_SLICE_X155Y123_CQ;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B3 = CLBLM_L_X98Y123_SLICE_X154Y123_AQ;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B4 = CLBLM_L_X98Y123_SLICE_X154Y123_A5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B5 = CLBLM_L_X98Y123_SLICE_X154Y123_C5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_T1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D3 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_D1 = CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C1 = CLBLM_L_X98Y123_SLICE_X155Y123_CQ;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C2 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C4 = CLBLM_R_X97Y122_SLICE_X152Y122_CQ;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C5 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_C6 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1 = 1'b0;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C3 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C4 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D1 = CLBLM_L_X98Y123_SLICE_X154Y123_C5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D2 = CLBLM_L_X98Y123_SLICE_X154Y123_AQ;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D3 = CLBLL_L_X102Y124_SLICE_X160Y124_D5Q;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D4 = CLBLM_L_X98Y123_SLICE_X155Y123_CQ;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_D6 = CLBLM_L_X98Y123_SLICE_X154Y123_A5Q;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1 = 1'b1;
  assign CLBLM_L_X98Y123_SLICE_X154Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y123_SLICE_X142Y123_D4 = 1'b1;
  assign LIOB33_X0Y63_IOB_X0Y64_O = 1'b0;
  assign LIOB33_X0Y63_IOB_X0Y63_O = 1'b0;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C4 = CLBLM_R_X97Y122_SLICE_X153Y122_DO6;
  assign LIOB33_X0Y63_IOB_X0Y64_T = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y63_IOB_X0Y63_T = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b0;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b0;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A1 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A2 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A3 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A4 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A5 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_A6 = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y151_T = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y152_T = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B1 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B2 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B3 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B4 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B5 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_B6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C1 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C2 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C3 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C4 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C5 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_C6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D1 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D2 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D3 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D4 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D5 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X151Y117_D6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A2 = CLBLM_R_X95Y118_SLICE_X150Y118_DO6;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A3 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A4 = CLBLM_L_X94Y117_SLICE_X149Y117_CO6;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A5 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_A6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B2 = CLBLM_R_X95Y117_SLICE_X150Y117_BQ;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B3 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B4 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B5 = CLBLM_R_X95Y117_SLICE_X150Y117_A5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_B6 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A1 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A2 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A3 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A4 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A5 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_A6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C1 = CLBLM_R_X95Y118_SLICE_X150Y118_C5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C2 = CLBLM_R_X95Y117_SLICE_X150Y117_CQ;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B1 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B2 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B3 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B4 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B5 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_B6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C1 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C2 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C3 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C4 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C5 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_C6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D2 = CLBLM_R_X95Y118_SLICE_X151Y118_A5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D3 = CLBLM_R_X95Y117_SLICE_X150Y117_BQ;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D4 = CLBLM_R_X95Y117_SLICE_X150Y117_A5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D5 = CLBLM_R_X95Y117_SLICE_X150Y117_B5Q;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_D6 = 1'b1;
  assign CLBLM_R_X95Y117_SLICE_X150Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D1 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D2 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D3 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D4 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D5 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X155Y124_D6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A2 = CLBLM_L_X98Y124_SLICE_X154Y124_B5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A3 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A4 = CLBLL_L_X100Y124_SLICE_X157Y124_BQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A5 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C1 = CLBLM_R_X93Y123_SLICE_X146Y123_BQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C2 = CLBLM_R_X93Y122_SLICE_X146Y122_A5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_A6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C3 = CLBLM_R_X97Y123_SLICE_X152Y123_CQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B2 = CLBLM_L_X98Y124_SLICE_X154Y124_BQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B3 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B4 = CLBLL_L_X100Y125_SLICE_X157Y125_CQ;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B5 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_B6 = 1'b1;
  assign CLBLM_R_X93Y123_SLICE_X146Y123_C5 = CLBLM_L_X92Y123_SLICE_X145Y123_CQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C1 = CLBLL_L_X100Y123_SLICE_X157Y123_AQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C2 = CLBLM_R_X97Y123_SLICE_X153Y123_DO6;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C3 = CLBLL_L_X100Y125_SLICE_X156Y125_CO6;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C4 = CLBLM_R_X97Y123_SLICE_X153Y123_A5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D2 = 1'b1;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D3 = CLBLM_L_X98Y124_SLICE_X154Y124_BQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D4 = CLBLM_L_X98Y124_SLICE_X154Y124_A5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D5 = CLBLM_L_X98Y124_SLICE_X154Y124_B5Q;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_D6 = CLBLL_L_X100Y125_SLICE_X157Y125_CQ;
  assign CLBLM_L_X98Y124_SLICE_X154Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y65_IOB_X0Y66_O = 1'b0;
  assign LIOB33_X0Y65_IOB_X0Y65_O = 1'b0;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = 1'b0;
  assign LIOB33_X0Y65_IOB_X0Y66_T = 1'b1;
  assign LIOB33_X0Y65_IOB_X0Y65_T = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y112_O = 1'b0;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b0;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b0;
  assign RIOB33_X105Y153_IOB_X1Y154_T = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_T = 1'b1;
  assign RIOB33_X105Y91_IOB_X1Y92_O = CLBLL_L_X102Y119_SLICE_X160Y119_CO6;
  assign RIOB33_X105Y91_IOB_X1Y91_O = CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_D1 = 1'b0;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A2 = CLBLM_R_X95Y117_SLICE_X150Y117_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A3 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A4 = CLBLM_R_X97Y119_SLICE_X152Y119_BQ;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A5 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_A6 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y112_T = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B2 = CLBLM_R_X95Y118_SLICE_X151Y118_BQ;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B3 = CLBLM_R_X95Y118_SLICE_X151Y118_AQ;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B4 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B5 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C1 = CLBLM_R_X97Y119_SLICE_X152Y119_BQ;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C3 = CLBLM_R_X95Y118_SLICE_X151Y118_BQ;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C4 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C5 = CLBLM_R_X95Y118_SLICE_X151Y118_AQ;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_C6 = CLBLM_R_X95Y118_SLICE_X151Y118_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D1 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D2 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D3 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D4 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D5 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_D6 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X95Y118_SLICE_X151Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A2 = CLBLM_R_X95Y118_SLICE_X151Y118_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A3 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A4 = CLBLM_R_X95Y118_SLICE_X150Y118_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A5 = CLBLM_L_X94Y118_SLICE_X148Y118_BO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_A6 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B2 = CLBLL_L_X100Y121_SLICE_X156Y121_C5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B3 = CLBLM_R_X95Y118_SLICE_X151Y118_A5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B4 = CLBLM_L_X94Y117_SLICE_X148Y117_CO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B5 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_B6 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A4 = CLBLM_L_X98Y125_SLICE_X155Y125_BO6;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A5 = CLBLM_L_X98Y126_SLICE_X154Y126_AQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_A6 = CLBLM_R_X103Y126_SLICE_X162Y126_DO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C1 = CLBLM_L_X98Y119_SLICE_X154Y119_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C2 = CLBLM_R_X95Y118_SLICE_X150Y118_CQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_AX = CLBLM_L_X98Y125_SLICE_X155Y125_BO5;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B2 = CLBLM_L_X98Y125_SLICE_X155Y125_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B3 = CLBLM_L_X98Y125_SLICE_X155Y125_AQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B4 = CLBLM_L_X98Y125_SLICE_X155Y125_CQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B5 = CLBLM_L_X98Y125_SLICE_X155Y125_C5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_B6 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C1 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C2 = CLBLM_L_X98Y125_SLICE_X155Y125_CQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C4 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C5 = CLBLM_L_X98Y125_SLICE_X155Y125_AQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_C6 = 1'b1;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D2 = CLBLL_L_X102Y121_SLICE_X161Y121_DO6;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D3 = CLBLM_R_X95Y117_SLICE_X150Y117_DO6;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D4 = CLBLM_R_X97Y119_SLICE_X152Y119_A5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D5 = CLBLM_R_X95Y118_SLICE_X150Y118_B5Q;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y118_SLICE_X150Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D1 = CLBLM_L_X98Y125_SLICE_X155Y125_C5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D3 = CLBLM_L_X98Y125_SLICE_X155Y125_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D4 = CLBLM_L_X98Y125_SLICE_X155Y125_AQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D5 = CLBLM_L_X98Y125_SLICE_X154Y125_DQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_D6 = CLBLM_L_X98Y125_SLICE_X155Y125_CQ;
  assign CLBLM_L_X98Y125_SLICE_X155Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A2 = CLBLM_L_X98Y127_SLICE_X155Y127_B5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A3 = CLBLM_R_X101Y126_SLICE_X159Y126_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A4 = CLBLM_L_X98Y128_SLICE_X154Y128_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A5 = CLBLM_R_X97Y124_SLICE_X153Y124_AO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_A6 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B2 = CLBLL_L_X100Y123_SLICE_X157Y123_AQ;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B3 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B4 = CLBLM_L_X98Y125_SLICE_X154Y125_B5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B5 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = 1'b0;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C1 = CLBLL_L_X100Y124_SLICE_X157Y124_B5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C2 = CLBLL_L_X100Y126_SLICE_X156Y126_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C4 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C5 = CLBLM_R_X97Y125_SLICE_X153Y125_CO6;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_C6 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D1 = CLBLM_R_X97Y126_SLICE_X153Y126_C5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D2 = CLBLM_R_X95Y125_SLICE_X150Y125_B5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D3 = CLBLM_L_X98Y125_SLICE_X154Y125_DQ;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D4 = CLBLM_R_X95Y124_SLICE_X151Y124_A5Q;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_D6 = 1'b1;
  assign CLBLM_L_X98Y125_SLICE_X154Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = 1'b0;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = 1'b0;
  assign LIOB33_X0Y67_IOB_X0Y68_O = 1'b0;
  assign LIOB33_X0Y67_IOB_X0Y67_O = 1'b0;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_D1 = 1'b0;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOB33_X0Y67_IOB_X0Y68_T = 1'b1;
  assign LIOB33_X0Y67_IOB_X0Y67_T = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_T1 = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_D1 = CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_D1 = 1'b0;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_D1 = 1'b0;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b0;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b0;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_D1 = CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y70_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_T = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_T = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_D1 = 1'b0;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_OLOGIC_X0Y69_T1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A1 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A2 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A3 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A4 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_A6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B1 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B2 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B3 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B4 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_B6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C1 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C2 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C3 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C4 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_C6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D1 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D2 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D3 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D4 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X151Y119_D6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A2 = CLBLM_R_X95Y119_SLICE_X150Y119_B5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A3 = CLBLM_R_X95Y118_SLICE_X150Y118_A5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A4 = CLBLM_L_X94Y119_SLICE_X149Y119_CO6;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_A6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B2 = CLBLM_R_X97Y120_SLICE_X153Y120_AQ;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B3 = CLBLM_R_X97Y119_SLICE_X153Y119_C5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B4 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B5 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_B6 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A3 = CLBLM_L_X98Y126_SLICE_X154Y126_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A4 = CLBLM_L_X98Y126_SLICE_X155Y126_BO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A5 = CLBLL_L_X102Y127_SLICE_X161Y127_DO6;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C2 = CLBLM_R_X95Y119_SLICE_X150Y119_CQ;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_C3 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_AX = CLBLM_L_X98Y126_SLICE_X155Y126_BO5;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B3 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B1 = CLBLM_L_X98Y126_SLICE_X155Y126_CQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B2 = CLBLM_L_X98Y126_SLICE_X155Y126_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B3 = CLBLM_L_X98Y126_SLICE_X155Y126_AQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B5 = CLBLM_L_X98Y126_SLICE_X155Y126_C5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_B6 = 1'b1;
  assign CLBLM_L_X94Y120_SLICE_X149Y120_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C1 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C2 = CLBLM_L_X98Y126_SLICE_X155Y126_CQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C4 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C5 = CLBLM_L_X98Y126_SLICE_X155Y126_AQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_C6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D1 = CLBLM_R_X95Y119_SLICE_X150Y119_C5Q;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D2 = CLBLM_R_X95Y119_SLICE_X150Y119_CQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D4 = CLBLM_R_X97Y120_SLICE_X153Y120_AQ;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_D6 = 1'b1;
  assign CLBLM_R_X95Y119_SLICE_X150Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D1 = CLBLM_L_X98Y126_SLICE_X155Y126_C5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D2 = CLBLM_L_X98Y126_SLICE_X155Y126_CQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D4 = CLBLM_L_X98Y126_SLICE_X155Y126_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D5 = CLBLM_L_X98Y126_SLICE_X155Y126_AQ;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_D6 = CLBLM_R_X97Y126_SLICE_X153Y126_C5Q;
  assign CLBLM_L_X98Y126_SLICE_X155Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A2 = CLBLM_L_X98Y126_SLICE_X154Y126_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A3 = CLBLM_R_X97Y129_SLICE_X152Y129_AQ;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A4 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A5 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_A6 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B2 = CLBLM_L_X98Y125_SLICE_X154Y125_C5Q;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B3 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B4 = CLBLL_L_X100Y126_SLICE_X156Y126_B5Q;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B5 = CLBLM_L_X98Y126_SLICE_X154Y126_CO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_B6 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C2 = CLBLL_L_X100Y127_SLICE_X156Y127_CO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C3 = CLBLM_R_X97Y125_SLICE_X153Y125_DO6;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C4 = CLBLM_R_X97Y125_SLICE_X152Y125_A5Q;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_C6 = CLBLM_L_X98Y125_SLICE_X154Y125_BQ;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D1 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D2 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D3 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D4 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D5 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_D6 = 1'b1;
  assign CLBLM_L_X98Y126_SLICE_X154Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y69_IOB_X0Y70_O = 1'b0;
  assign LIOB33_X0Y69_IOB_X0Y69_O = 1'b0;
  assign LIOB33_X0Y69_IOB_X0Y70_T = 1'b1;
  assign LIOB33_X0Y69_IOB_X0Y69_T = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A2 = CLBLM_R_X93Y122_SLICE_X146Y122_AQ;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b0;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b0;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A6 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_T = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y157_T = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B1 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B3 = CLBLM_R_X89Y120_SLICE_X140Y120_AQ;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C1 = CLBLM_R_X93Y121_SLICE_X146Y121_BQ;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C3 = CLBLM_R_X93Y122_SLICE_X147Y122_A5Q;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C4 = CLBLM_L_X92Y121_SLICE_X145Y121_C5Q;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C5 = CLBLM_L_X92Y121_SLICE_X144Y121_D5Q;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A1 = CLBLM_R_X97Y123_SLICE_X153Y123_AQ;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A2 = CLBLM_R_X95Y121_SLICE_X151Y121_B5Q;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A4 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A5 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_A6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B1 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B2 = CLBLM_R_X95Y120_SLICE_X151Y120_BQ;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B4 = CLBLM_R_X95Y120_SLICE_X151Y120_AQ;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B5 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_B6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C1 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C2 = CLBLM_R_X95Y120_SLICE_X151Y120_AQ;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C3 = CLBLM_R_X95Y120_SLICE_X151Y120_BQ;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C5 = CLBLM_R_X97Y123_SLICE_X153Y123_AQ;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_C6 = CLBLM_R_X95Y120_SLICE_X151Y120_B5Q;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D1 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D2 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D3 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D4 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D5 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_D6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X151Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A1 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A2 = CLBLM_R_X95Y120_SLICE_X150Y120_A5Q;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A3 = CLBLM_R_X95Y124_SLICE_X150Y124_AQ;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A4 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_A6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B1 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B2 = CLBLM_R_X95Y120_SLICE_X150Y120_BQ;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B3 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B4 = CLBLM_R_X95Y122_SLICE_X150Y122_BQ;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_B6 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A2 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A3 = CLBLM_L_X98Y127_SLICE_X154Y127_CO6;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A4 = CLBLM_L_X98Y127_SLICE_X154Y127_B5Q;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A5 = CLBLL_L_X100Y127_SLICE_X157Y127_B5Q;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_A6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C1 = CLBLM_R_X95Y122_SLICE_X150Y122_AQ;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C2 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B2 = CLBLM_L_X98Y127_SLICE_X155Y127_BQ;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B3 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B4 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B5 = CLBLM_L_X98Y128_SLICE_X154Y128_CQ;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_B6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D1 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C2 = CLBLM_L_X98Y128_SLICE_X154Y128_CQ;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C3 = CLBLM_L_X98Y127_SLICE_X155Y127_BQ;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C4 = CLBLM_R_X101Y128_SLICE_X158Y128_AQ;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C5 = CLBLM_L_X98Y127_SLICE_X155Y127_B5Q;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_C6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D2 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D3 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D4 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D5 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_D6 = 1'b1;
  assign CLBLM_R_X95Y120_SLICE_X150Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D1 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D2 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D3 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D4 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D5 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_D6 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X155Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A2 = CLBLM_L_X98Y127_SLICE_X154Y127_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A3 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A4 = CLBLM_L_X98Y125_SLICE_X154Y125_BQ;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A5 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_A6 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B2 = CLBLM_L_X98Y127_SLICE_X154Y127_DO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B3 = CLBLL_L_X100Y127_SLICE_X156Y127_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B4 = CLBLM_L_X98Y126_SLICE_X154Y126_B5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B5 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_B6 = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C2 = CLBLM_L_X98Y127_SLICE_X154Y127_AQ;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C3 = CLBLM_R_X101Y129_SLICE_X158Y129_DO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C4 = CLBLM_R_X97Y127_SLICE_X152Y127_DO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C5 = CLBLM_R_X97Y127_SLICE_X153Y127_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y71_IOB_X0Y71_O = 1'b0;
  assign LIOB33_X0Y71_IOB_X0Y72_O = 1'b0;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y71_IOB_X0Y72_T = 1'b1;
  assign LIOB33_X0Y71_IOB_X0Y71_T = 1'b1;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D2 = CLBLM_R_X97Y126_SLICE_X152Y126_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D3 = CLBLL_L_X100Y127_SLICE_X157Y127_CO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D4 = CLBLM_L_X98Y127_SLICE_X154Y127_A5Q;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D5 = CLBLM_R_X97Y126_SLICE_X152Y126_CO6;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y124_SLICE_X143Y124_C2 = CLBLM_L_X90Y124_SLICE_X143Y124_CQ;
  assign CLBLM_L_X98Y127_SLICE_X154Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y159_IOB_X1Y160_O = 1'b0;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b0;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B4 = CLBLM_L_X90Y122_SLICE_X142Y122_BQ;
  assign RIOB33_X105Y159_IOB_X1Y160_T = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y159_T = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = 1'b0;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C2 = CLBLM_L_X92Y122_SLICE_X144Y122_CQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C3 = CLBLM_L_X90Y120_SLICE_X142Y120_B5Q;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D2 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = 1'b0;
  assign LIOI3_TBYTETERM_X0Y213_OLOGIC_X0Y214_D1 = 1'b0;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = 1'b0;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A1 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A2 = CLBLM_R_X97Y121_SLICE_X152Y121_BQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A4 = CLBLM_R_X95Y121_SLICE_X151Y121_AQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A5 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_A6 = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_D1 = 1'b0;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B1 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B2 = CLBLM_R_X95Y121_SLICE_X151Y121_BQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B4 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B5 = CLBLM_R_X97Y121_SLICE_X153Y121_BQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_B6 = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_T1 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_D1 = 1'b0;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C1 = CLBLM_R_X97Y121_SLICE_X152Y121_AQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C2 = CLBLM_R_X97Y121_SLICE_X152Y121_BQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C3 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C4 = CLBLM_R_X95Y121_SLICE_X151Y121_A5Q;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_C6 = CLBLM_R_X95Y121_SLICE_X151Y121_AQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_D1 = 1'b0;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_T1 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D1 = CLBLM_R_X95Y121_SLICE_X151Y121_BQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D3 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D4 = CLBLM_R_X97Y121_SLICE_X153Y121_BQ;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D5 = CLBLM_R_X95Y121_SLICE_X151Y121_B5Q;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_D6 = CLBLM_R_X95Y120_SLICE_X151Y120_A5Q;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_D1 = 1'b0;
  assign CLBLM_R_X95Y121_SLICE_X151Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y82_T1 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A1 = CLBLM_R_X97Y121_SLICE_X152Y121_B5Q;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A6 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A2 = CLBLM_L_X94Y120_SLICE_X148Y120_B5Q;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A4 = CLBLM_R_X95Y121_SLICE_X151Y121_A5Q;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A5 = CLBLM_R_X95Y121_SLICE_X150Y121_AQ;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_A6 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1 = 1'b0;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B3 = CLBLM_R_X95Y121_SLICE_X151Y121_CO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B4 = CLBLM_R_X101Y121_SLICE_X158Y121_CO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B5 = CLBLM_R_X95Y120_SLICE_X150Y120_AQ;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_B6 = CLBLM_R_X95Y121_SLICE_X150Y121_A5Q;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_D1 = 1'b0;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A1 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A2 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A3 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A4 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A5 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_A6 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C1 = CLBLM_R_X95Y120_SLICE_X150Y120_A5Q;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C2 = CLBLM_R_X95Y121_SLICE_X150Y121_AQ;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_C3 = CLBLM_R_X97Y121_SLICE_X152Y121_DO6;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B1 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B2 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B3 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B4 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B5 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_B6 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D1 = CLBLM_R_X95Y124_SLICE_X150Y124_AQ;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D2 = CLBLM_L_X94Y120_SLICE_X148Y120_B5Q;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C1 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C2 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C3 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C4 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C5 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_C6 = 1'b1;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D3 = CLBLM_L_X98Y122_SLICE_X155Y122_DO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D4 = CLBLM_R_X95Y120_SLICE_X150Y120_CO6;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y121_SLICE_X150Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D1 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D2 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D3 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D4 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D5 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X155Y128_D6 = 1'b1;
  assign LIOB33_X0Y73_IOB_X0Y73_O = 1'b0;
  assign LIOB33_X0Y73_IOB_X0Y74_O = 1'b0;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A2 = CLBLM_L_X98Y128_SLICE_X154Y128_C5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A3 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A4 = CLBLM_R_X97Y124_SLICE_X152Y124_CO6;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A5 = CLBLM_R_X97Y127_SLICE_X153Y127_A5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_A6 = 1'b1;
  assign LIOB33_X0Y73_IOB_X0Y73_T = 1'b1;
  assign LIOB33_X0Y73_IOB_X0Y74_T = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B2 = CLBLM_L_X98Y128_SLICE_X154Y128_BQ;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B3 = CLBLL_L_X100Y129_SLICE_X157Y129_AQ;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B4 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B5 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_B6 = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_T1 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C1 = CLBLM_R_X101Y128_SLICE_X158Y128_AQ;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C2 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C3 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C5 = CLBLM_L_X98Y128_SLICE_X154Y128_B5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_C6 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y161_IOB_X1Y161_O = 1'b0;
  assign RIOB33_X105Y161_IOB_X1Y162_O = 1'b0;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D1 = CLBLM_L_X98Y128_SLICE_X154Y128_C5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D2 = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D3 = CLBLM_L_X98Y128_SLICE_X154Y128_BQ;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D4 = CLBLL_L_X100Y129_SLICE_X157Y129_AQ;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D5 = CLBLM_L_X98Y128_SLICE_X154Y128_B5Q;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOB33_X105Y161_IOB_X1Y161_T = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_T = 1'b1;
  assign CLBLM_L_X98Y128_SLICE_X154Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y124_SLICE_X142Y124_D1 = CLBLM_L_X90Y124_SLICE_X142Y124_C5Q;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_T1 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C4 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C5 = CLBLM_R_X95Y124_SLICE_X150Y124_BQ;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C6 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A1 = CLBLM_R_X97Y125_SLICE_X152Y125_CO6;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A2 = CLBLM_L_X94Y120_SLICE_X149Y120_A5Q;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A4 = CLBLM_R_X97Y121_SLICE_X153Y121_AQ;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_A6 = CLBLM_R_X95Y120_SLICE_X151Y120_CO6;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B1 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B2 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B3 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B4 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B5 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_B6 = 1'b1;
  assign CLBLM_R_X101Y135_SLICE_X158Y135_D5 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C1 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C2 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C3 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C4 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C5 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_C6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B4 = CLBLM_L_X94Y125_SLICE_X149Y125_DQ;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D1 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D2 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D3 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D4 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D5 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X151Y122_D6 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D3 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A1 = CLBLM_R_X95Y124_SLICE_X150Y124_B5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A2 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A4 = CLBLM_R_X95Y121_SLICE_X150Y121_DO6;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A5 = CLBLM_R_X97Y123_SLICE_X152Y123_B5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_A6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B5 = CLBLM_L_X94Y125_SLICE_X149Y125_C5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B1 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D3 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B2 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B4 = CLBLM_R_X95Y122_SLICE_X150Y122_AQ;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B5 = CLBLM_R_X95Y122_SLICE_X150Y122_C5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_B6 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A1 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A2 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A3 = CLBLM_L_X98Y129_SLICE_X155Y129_AQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A5 = CLBLM_L_X98Y127_SLICE_X154Y127_AQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_A6 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C2 = CLBLM_R_X95Y122_SLICE_X150Y122_CQ;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_C3 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B1 = CLBLM_L_X98Y129_SLICE_X154Y129_AQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B2 = CLBLM_L_X98Y130_SLICE_X155Y130_BQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B3 = CLBLM_L_X98Y129_SLICE_X155Y129_CQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B5 = CLBLM_L_X98Y129_SLICE_X155Y129_C5Q;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_B6 = 1'b1;
  assign CLBLM_L_X94Y125_SLICE_X149Y125_B6 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C1 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C3 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C4 = CLBLM_L_X98Y130_SLICE_X155Y130_BQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C5 = CLBLM_L_X98Y129_SLICE_X155Y129_CQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_C6 = 1'b1;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D1 = CLBLM_R_X95Y122_SLICE_X150Y122_C5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D2 = CLBLM_R_X95Y122_SLICE_X150Y122_CQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D5 = CLBLM_R_X95Y122_SLICE_X150Y122_B5Q;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_D6 = CLBLM_R_X95Y124_SLICE_X150Y124_BQ;
  assign CLBLM_R_X95Y122_SLICE_X150Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D1 = CLBLM_L_X98Y129_SLICE_X155Y129_C5Q;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D3 = CLBLM_L_X98Y130_SLICE_X155Y130_BQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D4 = CLBLM_R_X97Y130_SLICE_X153Y130_AQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D5 = CLBLM_L_X98Y129_SLICE_X154Y129_AQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_D6 = CLBLM_L_X98Y129_SLICE_X155Y129_CQ;
  assign CLBLM_L_X98Y129_SLICE_X155Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y113_IOB_X0Y114_O = 1'b0;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A1 = CLBLM_L_X98Y129_SLICE_X154Y129_B5Q;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A3 = CLBLM_L_X98Y129_SLICE_X154Y129_CQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A4 = CLBLM_L_X98Y130_SLICE_X155Y130_CQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A5 = CLBLM_L_X98Y129_SLICE_X154Y129_BQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_A6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y113_O = 1'b0;
  assign RIOB33_X105Y163_IOB_X1Y163_O = 1'b0;
  assign RIOB33_X105Y163_IOB_X1Y164_O = 1'b0;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_AX = CLBLM_L_X98Y129_SLICE_X155Y129_BO5;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B2 = CLBLM_L_X98Y129_SLICE_X154Y129_BQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B3 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B4 = CLBLM_L_X98Y130_SLICE_X155Y130_CQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B5 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_B6 = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y163_T = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y164_T = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C1 = CLBLM_L_X98Y129_SLICE_X154Y129_BQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C2 = CLBLM_L_X98Y129_SLICE_X154Y129_CQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C3 = CLBLM_R_X97Y129_SLICE_X152Y129_BQ;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C5 = CLBLM_L_X98Y129_SLICE_X154Y129_B5Q;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_C6 = CLBLM_L_X98Y130_SLICE_X155Y130_CQ;
  assign RIOB33_X105Y93_IOB_X1Y93_O = CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  assign RIOB33_X105Y93_IOB_X1Y94_O = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_CX = CLBLM_L_X98Y129_SLICE_X154Y129_AO5;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D1 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D2 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D3 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D4 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D5 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_D6 = 1'b1;
  assign CLBLM_L_X98Y129_SLICE_X154Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y113_IOB_X0Y114_T = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y113_T = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A1 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A3 = CLBLM_R_X97Y121_SLICE_X153Y121_AQ;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A4 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A5 = CLBLM_R_X95Y123_SLICE_X151Y123_A5Q;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_A6 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B1 = CLBLM_R_X95Y123_SLICE_X151Y123_BQ;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B3 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B4 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B5 = CLBLM_R_X95Y123_SLICE_X150Y123_AQ;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_B6 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C1 = CLBLM_L_X94Y122_SLICE_X149Y122_B5Q;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C2 = CLBLM_R_X95Y123_SLICE_X150Y123_CO6;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C4 = CLBLM_R_X95Y123_SLICE_X151Y123_A5Q;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C5 = CLBLM_R_X97Y125_SLICE_X153Y125_DO6;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D1 = CLBLM_R_X95Y123_SLICE_X150Y123_AQ;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D2 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D3 = CLBLM_R_X97Y125_SLICE_X152Y125_AQ;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D4 = CLBLM_R_X95Y123_SLICE_X151Y123_BQ;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D5 = CLBLM_R_X95Y123_SLICE_X151Y123_B5Q;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y123_SLICE_X151Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y77_IOB_X0Y78_O = 1'b0;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A1 = CLBLM_R_X95Y123_SLICE_X150Y123_B5Q;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A2 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A3 = CLBLM_R_X97Y125_SLICE_X152Y125_AQ;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A5 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_A6 = 1'b1;
  assign LIOB33_X0Y77_IOB_X0Y77_O = 1'b0;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B1 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B2 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B3 = CLBLM_R_X97Y123_SLICE_X152Y123_AQ;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B5 = CLBLM_R_X95Y123_SLICE_X150Y123_BQ;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_B6 = 1'b1;
  assign LIOB33_X0Y77_IOB_X0Y77_T = 1'b1;
  assign LIOB33_X0Y77_IOB_X0Y78_T = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A1 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A2 = CLBLM_L_X98Y130_SLICE_X155Y130_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A3 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A5 = CLBLM_L_X98Y129_SLICE_X155Y129_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_A6 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C1 = CLBLM_R_X95Y123_SLICE_X150Y123_BQ;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C2 = CLBLM_R_X97Y123_SLICE_X152Y123_AQ;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C3 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B1 = CLBLM_R_X101Y130_SLICE_X159Y130_DO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B4 = CLBLM_L_X98Y129_SLICE_X155Y129_BO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B5 = CLBLM_L_X98Y130_SLICE_X155Y130_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D1 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C1 = CLBLM_L_X98Y129_SLICE_X154Y129_AO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C4 = CLBLL_L_X102Y131_SLICE_X160Y131_DO6;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_C6 = CLBLM_L_X98Y129_SLICE_X155Y129_A5Q;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D6 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D5 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y165_T = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y166_T = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D1 = CLBLM_L_X98Y128_SLICE_X154Y128_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D3 = CLBLM_L_X98Y132_SLICE_X155Y132_CQ;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D4 = CLBLM_L_X98Y129_SLICE_X154Y129_CQ;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D5 = CLBLM_R_X97Y130_SLICE_X152Y130_AQ;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_D6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = 1'b0;
  assign CLBLM_L_X98Y130_SLICE_X155Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A1 = CLBLL_L_X102Y130_SLICE_X160Y130_DO6;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A3 = CLBLM_L_X98Y133_SLICE_X154Y133_AQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A4 = CLBLM_L_X98Y130_SLICE_X154Y130_BO6;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_D1 = 1'b0;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_AX = CLBLM_L_X98Y130_SLICE_X154Y130_BO5;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B2 = CLBLM_L_X98Y130_SLICE_X154Y130_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B3 = CLBLM_L_X98Y130_SLICE_X154Y130_AQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B4 = CLBLM_L_X98Y130_SLICE_X154Y130_CQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B5 = CLBLM_L_X98Y130_SLICE_X154Y130_C5Q;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_B6 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_T1 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_D1 = 1'b0;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C1 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C2 = CLBLM_L_X98Y130_SLICE_X154Y130_CQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C3 = CLBLM_L_X98Y130_SLICE_X154Y130_AQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C5 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_C6 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_D1 = 1'b0;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_T1 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_D1 = 1'b0;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_T1 = 1'b1;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D1 = CLBLM_L_X98Y130_SLICE_X154Y130_C5Q;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D2 = CLBLM_L_X98Y130_SLICE_X154Y130_AQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D4 = CLBLM_L_X98Y130_SLICE_X154Y130_A5Q;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D5 = CLBLM_L_X98Y130_SLICE_X154Y130_CQ;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_D6 = CLBLM_R_X97Y129_SLICE_X152Y129_CQ;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_T1 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_D1 = 1'b0;
  assign CLBLM_L_X98Y130_SLICE_X154Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1 = CLBLM_R_X101Y117_SLICE_X159Y117_AO5;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_D1 = 1'b0;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1 = CLBLL_L_X100Y115_SLICE_X157Y115_CO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A1 = CLBLL_L_X100Y124_SLICE_X156Y124_CO6;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A3 = CLBLM_R_X95Y124_SLICE_X151Y124_BO6;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A5 = CLBLM_R_X95Y125_SLICE_X150Y125_AQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_AX = CLBLM_R_X95Y124_SLICE_X151Y124_BO5;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B1 = CLBLM_R_X95Y124_SLICE_X151Y124_CQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B3 = CLBLM_R_X95Y124_SLICE_X151Y124_AQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B4 = CLBLM_R_X97Y124_SLICE_X152Y124_B5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B5 = CLBLM_R_X95Y124_SLICE_X151Y124_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_B6 = 1'b1;
  assign LIOB33_X0Y79_IOB_X0Y80_O = 1'b0;
  assign LIOB33_X0Y79_IOB_X0Y79_O = 1'b0;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C1 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C2 = CLBLM_L_X94Y125_SLICE_X149Y125_CQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C3 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C5 = CLBLM_R_X95Y124_SLICE_X151Y124_AQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_C6 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y79_IOB_X0Y79_T = 1'b1;
  assign LIOB33_X0Y79_IOB_X0Y80_T = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D1 = CLBLM_L_X94Y124_SLICE_X148Y124_C5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D2 = CLBLM_R_X95Y124_SLICE_X151Y124_CQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D4 = CLBLM_R_X95Y124_SLICE_X151Y124_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D5 = CLBLM_R_X95Y124_SLICE_X151Y124_AQ;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_D6 = CLBLM_R_X97Y124_SLICE_X152Y124_B5Q;
  assign CLBLM_R_X95Y124_SLICE_X151Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A1 = CLBLM_L_X94Y124_SLICE_X148Y124_AQ;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A2 = CLBLM_R_X95Y124_SLICE_X150Y124_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A3 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A5 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_A6 = 1'b1;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_D1 = 1'b0;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = 1'b0;
  assign RIOB33_X105Y167_IOB_X1Y168_O = 1'b0;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B1 = CLBLM_R_X95Y124_SLICE_X150Y124_DO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B2 = CLBLM_L_X98Y125_SLICE_X154Y125_D5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B3 = CLBLM_L_X94Y128_SLICE_X149Y128_C5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B5 = CLBLM_R_X95Y124_SLICE_X150Y124_C5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_B6 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y168_T = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A2 = CLBLM_L_X98Y131_SLICE_X155Y131_A5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A3 = CLBLM_L_X98Y130_SLICE_X155Y130_AQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A6 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C1 = CLBLM_L_X94Y124_SLICE_X149Y124_BO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C2 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C3 = CLBLM_L_X94Y125_SLICE_X148Y125_B5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B1 = CLBLM_R_X97Y130_SLICE_X152Y130_AO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B3 = CLBLM_L_X98Y131_SLICE_X155Y131_AQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B4 = CLBLM_R_X101Y132_SLICE_X159Y132_DO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_BX = CLBLM_L_X98Y131_SLICE_X155Y131_CO5;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C1 = CLBLM_R_X97Y131_SLICE_X153Y131_BQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C2 = CLBLM_R_X97Y131_SLICE_X153Y131_B5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C4 = CLBLM_L_X98Y132_SLICE_X155Y132_BQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C5 = CLBLM_L_X98Y131_SLICE_X155Y131_B5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C6 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D2 = CLBLM_R_X97Y123_SLICE_X152Y123_DO6;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D3 = CLBLM_R_X95Y122_SLICE_X150Y122_DO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D4 = CLBLM_R_X95Y124_SLICE_X150Y124_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D5 = CLBLM_L_X94Y120_SLICE_X148Y120_C5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D2 = CLBLM_L_X98Y131_SLICE_X154Y131_A5Q;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D3 = CLBLM_L_X98Y131_SLICE_X155Y131_DQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D4 = CLBLM_L_X98Y129_SLICE_X154Y129_AQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D5 = CLBLM_L_X98Y130_SLICE_X155Y130_DQ;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D6 = 1'b1;
  assign LIOI3_X0Y75_OLOGIC_X0Y76_T1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = 1'b0;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A3 = CLBLM_R_X101Y131_SLICE_X158Y131_DO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A4 = CLBLM_L_X98Y131_SLICE_X154Y131_BO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A5 = CLBLM_L_X98Y130_SLICE_X155Y130_AQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_AX = CLBLM_L_X98Y131_SLICE_X154Y131_BO5;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B2 = CLBLM_L_X98Y131_SLICE_X154Y131_A5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B3 = CLBLM_L_X98Y131_SLICE_X154Y131_AQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B4 = CLBLM_L_X98Y131_SLICE_X154Y131_CQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B5 = CLBLM_L_X98Y131_SLICE_X154Y131_C5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C2 = CLBLM_L_X98Y131_SLICE_X154Y131_CQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C3 = CLBLM_L_X98Y131_SLICE_X154Y131_AQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C6 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C4 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A2 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A4 = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A5 = CLBLL_L_X102Y111_SLICE_X161Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D1 = CLBLM_L_X98Y131_SLICE_X154Y131_C5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D4 = CLBLM_L_X98Y131_SLICE_X154Y131_A5Q;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D6 = CLBLM_R_X97Y130_SLICE_X153Y130_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B2 = CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B3 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B4 = CLBLM_R_X101Y112_SLICE_X158Y112_BQ;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B5 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B6 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C1 = CLBLL_L_X102Y111_SLICE_X161Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C3 = CLBLL_L_X102Y111_SLICE_X161Y111_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C4 = CLBLM_R_X101Y112_SLICE_X158Y112_CO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C5 = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_D1 = 1'b0;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D2 = CLBLM_R_X101Y112_SLICE_X159Y112_C5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D3 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D4 = CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D5 = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D6 = CLBLM_R_X101Y112_SLICE_X158Y112_BQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A1 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A2 = CLBLM_L_X92Y123_SLICE_X145Y123_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A4 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A3 = CLBLL_L_X102Y111_SLICE_X161Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A4 = CLBLM_R_X103Y112_SLICE_X162Y112_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A5 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A6 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A5 = CLBLM_L_X92Y123_SLICE_X144Y123_AQ;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_A6 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B2 = CLBLL_L_X102Y111_SLICE_X161Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B3 = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B4 = CLBLM_R_X101Y112_SLICE_X159Y112_C5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B5 = CLBLM_R_X103Y112_SLICE_X162Y112_C5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B6 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D6 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C1 = CLBLL_L_X102Y111_SLICE_X161Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C3 = CLBLM_R_X103Y112_SLICE_X162Y112_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C5 = CLBLL_L_X100Y111_SLICE_X156Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C6 = CLBLL_L_X102Y111_SLICE_X161Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_CX = CLBLM_R_X103Y111_SLICE_X162Y111_AO5;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D1 = CLBLM_R_X103Y111_SLICE_X162Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D2 = CLBLM_R_X101Y111_SLICE_X158Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D3 = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D6 = CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y81_IOB_X0Y82_O = 1'b0;
  assign LIOB33_X0Y81_IOB_X0Y81_O = 1'b0;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOB33_X0Y81_IOB_X0Y82_T = 1'b1;
  assign LIOB33_X0Y81_IOB_X0Y81_T = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A1 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A2 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A4 = CLBLM_R_X95Y125_SLICE_X151Y125_AQ;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A5 = CLBLM_R_X95Y126_SLICE_X150Y126_AQ;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_A6 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B1 = CLBLM_R_X95Y123_SLICE_X151Y123_DO6;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B2 = CLBLM_R_X97Y126_SLICE_X152Y126_CO6;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B3 = CLBLM_R_X95Y123_SLICE_X151Y123_AQ;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B4 = CLBLM_L_X94Y122_SLICE_X149Y122_A5Q;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C1 = CLBLM_R_X95Y126_SLICE_X150Y126_AQ;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C2 = CLBLM_R_X97Y127_SLICE_X153Y127_AQ;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C4 = CLBLM_R_X95Y125_SLICE_X151Y125_A5Q;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C5 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_C6 = CLBLM_R_X95Y125_SLICE_X151Y125_AQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = 1'b0;
  assign RIOB33_X105Y169_IOB_X1Y170_O = 1'b0;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D1 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D2 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D3 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D4 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D5 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_D6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_T = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_T = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X151Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A1 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A2 = CLBLM_R_X95Y125_SLICE_X150Y125_A5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A4 = CLBLM_L_X94Y127_SLICE_X149Y127_AQ;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A5 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_A6 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B2 = CLBLM_R_X95Y125_SLICE_X150Y125_A5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B4 = CLBLM_L_X98Y125_SLICE_X155Y125_DO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_B6 = CLBLM_R_X95Y125_SLICE_X150Y125_CO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_BX = CLBLM_R_X95Y125_SLICE_X150Y125_CO5;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A1 = CLBLM_L_X98Y133_SLICE_X155Y133_BQ;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A2 = CLBLM_R_X97Y132_SLICE_X153Y132_AQ;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A4 = CLBLM_R_X97Y132_SLICE_X153Y132_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A5 = CLBLM_L_X98Y132_SLICE_X155Y132_AQ;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A6 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C2 = CLBLM_R_X95Y125_SLICE_X150Y125_B5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C3 = CLBLM_R_X95Y125_SLICE_X150Y125_BQ;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B1 = CLBLM_L_X98Y131_SLICE_X155Y131_CO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B4 = CLBLM_R_X101Y133_SLICE_X158Y133_DO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B5 = CLBLM_L_X98Y131_SLICE_X155Y131_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C4 = CLBLL_L_X102Y131_SLICE_X160Y131_BQ;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C1 = CLBLM_L_X98Y130_SLICE_X155Y130_D5Q;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C3 = CLBLM_L_X98Y131_SLICE_X155Y131_B5Q;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C4 = CLBLM_L_X98Y131_SLICE_X155Y131_D5Q;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C5 = CLBLM_L_X98Y132_SLICE_X155Y132_AQ;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C6 = 1'b1;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D1 = CLBLM_R_X95Y124_SLICE_X151Y124_C5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D4 = CLBLM_L_X94Y125_SLICE_X149Y125_CQ;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D5 = CLBLM_R_X95Y125_SLICE_X150Y125_B5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D6 = CLBLM_L_X94Y124_SLICE_X148Y124_CQ;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D5 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A1 = CLBLM_R_X93Y112_SLICE_X146Y112_B5Q;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A5 = CLBLM_R_X93Y115_SLICE_X146Y115_AQ;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_A6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B1 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B3 = CLBLM_L_X92Y112_SLICE_X145Y112_AQ;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B4 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B5 = CLBLM_L_X92Y112_SLICE_X145Y112_BQ;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_B6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A2 = CLBLM_L_X98Y133_SLICE_X154Y133_BQ;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A3 = CLBLM_R_X101Y133_SLICE_X159Y133_BO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A4 = CLBLM_L_X98Y132_SLICE_X154Y132_BO6;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C2 = CLBLM_L_X92Y112_SLICE_X145Y112_AQ;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C4 = CLBLM_L_X92Y112_SLICE_X145Y112_BQ;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C5 = CLBLM_L_X92Y112_SLICE_X145Y112_B5Q;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_C6 = CLBLM_R_X93Y115_SLICE_X146Y115_AQ;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_AX = CLBLM_L_X98Y132_SLICE_X154Y132_BO5;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B2 = CLBLM_L_X98Y132_SLICE_X154Y132_A5Q;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B3 = CLBLM_L_X98Y132_SLICE_X154Y132_AQ;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B4 = CLBLM_L_X98Y132_SLICE_X154Y132_CQ;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B5 = CLBLM_L_X98Y132_SLICE_X154Y132_C5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D1 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D2 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D4 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D5 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_D6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A3 = CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  assign CLBLM_L_X92Y112_SLICE_X145Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A4 = CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A5 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B2 = CLBLM_R_X101Y112_SLICE_X159Y112_CQ;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A1 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A2 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A4 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A5 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_A6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B4 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B5 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B6 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B1 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B2 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B4 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B5 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_B6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C4 = CLBLL_L_X100Y112_SLICE_X156Y112_CO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_CX = CLBLL_L_X102Y111_SLICE_X160Y111_AO5;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C1 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C2 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C4 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C5 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_C6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D1 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D2 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D3 = CLBLL_L_X100Y112_SLICE_X157Y112_AQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D4 = CLBLM_R_X101Y112_SLICE_X159Y112_CQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D5 = CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D1 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D2 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D3 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D4 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D5 = 1'b1;
  assign CLBLM_L_X92Y112_SLICE_X144Y112_D6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = 1'b0;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A2 = CLBLL_L_X102Y113_SLICE_X161Y113_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A3 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A4 = CLBLM_R_X101Y110_SLICE_X158Y110_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A5 = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B2 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B3 = CLBLL_L_X102Y113_SLICE_X161Y113_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B4 = CLBLM_R_X103Y112_SLICE_X163Y112_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B5 = CLBLM_R_X103Y112_SLICE_X162Y112_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = 1'b0;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_D1 = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C1 = CLBLM_R_X103Y112_SLICE_X163Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C2 = CLBLM_R_X103Y112_SLICE_X163Y112_BO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C4 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C6 = CLBLM_R_X101Y110_SLICE_X158Y110_CO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_T1 = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_D1 = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D2 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D3 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D4 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D5 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D6 = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_D1 = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = 1'b0;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_T1 = 1'b1;
  assign LIOB33_X0Y83_IOB_X0Y84_O = 1'b0;
  assign LIOB33_X0Y83_IOB_X0Y83_O = 1'b0;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOB33_X0Y83_IOB_X0Y84_T = 1'b1;
  assign LIOB33_X0Y83_IOB_X0Y83_T = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A2 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y171_O = 1'b0;
  assign RIOB33_X105Y171_IOB_X1Y172_O = 1'b0;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A2 = CLBLM_R_X95Y126_SLICE_X151Y126_A5Q;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A3 = CLBLM_R_X95Y123_SLICE_X151Y123_AQ;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_A6 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y171_T = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_T = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B1 = CLBLM_R_X97Y127_SLICE_X152Y127_DO6;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A2 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B4 = CLBLM_R_X95Y126_SLICE_X150Y126_CO6;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B5 = CLBLM_L_X94Y125_SLICE_X148Y125_B5Q;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_B6 = CLBLM_R_X95Y126_SLICE_X151Y126_A5Q;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A3 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C2 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C3 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A4 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C4 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_C6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_A6 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D2 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D3 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D4 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_D6 = 1'b1;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y126_SLICE_X151Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_B2 = CLBLM_L_X90Y123_SLICE_X142Y123_BQ;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A1 = CLBLM_R_X95Y126_SLICE_X150Y126_B5Q;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A2 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A3 = CLBLM_R_X97Y127_SLICE_X153Y127_AQ;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_A6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B1 = CLBLM_R_X95Y126_SLICE_X150Y126_BQ;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B3 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B4 = CLBLM_R_X97Y126_SLICE_X152Y126_AQ;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B2 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_B6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B3 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A2 = CLBLM_L_X98Y133_SLICE_X155Y133_A5Q;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A3 = CLBLM_L_X98Y131_SLICE_X155Y131_AQ;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A4 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A5 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_A6 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B2 = CLBLM_L_X98Y133_SLICE_X155Y133_A5Q;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B4 = CLBLL_L_X100Y134_SLICE_X156Y134_CO6;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B5 = CLBLM_L_X98Y132_SLICE_X155Y132_AO6;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B6 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C1 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C2 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C3 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C5 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_C6 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D1 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D2 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D4 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D5 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_D6 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D1 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D2 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D3 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D4 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D5 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_D6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C1 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A1 = CLBLM_R_X93Y114_SLICE_X146Y114_CO6;
  assign CLBLM_L_X98Y133_SLICE_X155Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A2 = CLBLM_R_X93Y113_SLICE_X146Y113_A5Q;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A3 = CLBLM_L_X92Y112_SLICE_X145Y112_B5Q;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C2 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_A5 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_A4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B1 = CLBLM_L_X92Y113_SLICE_X145Y113_B5Q;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B2 = CLBLM_L_X94Y113_SLICE_X148Y113_BQ;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B3 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C3 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_B4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C1 = CLBLM_L_X92Y113_SLICE_X145Y113_BQ;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C2 = CLBLM_L_X94Y116_SLICE_X148Y116_CO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C4 = CLBLM_L_X92Y113_SLICE_X145Y113_A5Q;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_C6 = CLBLM_L_X92Y112_SLICE_X145Y112_CO6;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A1 = CLBLL_L_X102Y111_SLICE_X161Y111_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A2 = CLBLM_R_X101Y113_SLICE_X158Y113_A5Q;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A3 = CLBLL_L_X102Y113_SLICE_X160Y113_AQ;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A4 = CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D2 = CLBLM_R_X93Y118_SLICE_X147Y118_CO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y113_SLICE_X145Y113_D5 = CLBLM_L_X92Y113_SLICE_X145Y113_B5Q;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C1 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_D5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C5 = 1'b1;
  assign CLBLM_L_X98Y133_SLICE_X154Y133_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A5 = CLBLM_L_X92Y113_SLICE_X145Y113_AQ;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_A6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C1 = CLBLM_L_X92Y113_SLICE_X145Y113_AQ;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C2 = CLBLM_L_X92Y113_SLICE_X144Y113_AQ;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C3 = CLBLM_L_X92Y113_SLICE_X144Y113_BQ;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C5 = CLBLM_L_X92Y113_SLICE_X144Y113_B5Q;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_C6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D6 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_D3 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D1 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D2 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D3 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D5 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_D6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D4 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D4 = 1'b1;
  assign CLBLM_L_X92Y113_SLICE_X144Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A2 = CLBLM_R_X101Y112_SLICE_X159Y112_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A3 = CLBLL_L_X102Y114_SLICE_X160Y114_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A5 = CLBLL_L_X102Y113_SLICE_X161Y113_CO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B2 = CLBLL_L_X102Y113_SLICE_X161Y113_BQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B3 = CLBLL_L_X102Y114_SLICE_X161Y114_A5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B4 = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B5 = CLBLL_L_X102Y115_SLICE_X161Y115_C5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C1 = CLBLM_R_X101Y112_SLICE_X159Y112_DO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C2 = CLBLM_R_X103Y113_SLICE_X162Y113_CO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C5 = CLBLL_L_X102Y113_SLICE_X161Y113_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C6 = CLBLM_R_X103Y113_SLICE_X163Y113_AQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y85_IOB_X0Y86_O = 1'b0;
  assign LIOB33_X0Y85_IOB_X0Y85_O = 1'b0;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D1 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D2 = CLBLM_R_X101Y113_SLICE_X159Y113_DO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D4 = CLBLL_L_X102Y113_SLICE_X161Y113_BQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D6 = CLBLL_L_X102Y114_SLICE_X161Y114_BO6;
  assign LIOB33_X0Y85_IOB_X0Y86_T = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y85_IOB_X0Y85_T = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = 1'b0;
  assign RIOB33_X105Y173_IOB_X1Y173_O = 1'b0;
  assign LIOB33_X0Y115_IOB_X0Y116_O = 1'b0;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b0;
  assign LIOB33_X0Y115_IOB_X0Y115_O = 1'b0;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A4 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y173_T = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_T = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C4 = CLBLM_R_X95Y123_SLICE_X150Y123_A5Q;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C5 = CLBLM_R_X95Y123_SLICE_X150Y123_B5Q;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOB33_X105Y95_IOB_X1Y96_O = CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  assign RIOB33_X105Y95_IOB_X1Y95_O = CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B2 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y116_T = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B5 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y115_T = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B6 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D2 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D3 = 1'b1;
  assign CLBLM_R_X95Y123_SLICE_X150Y123_D4 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A1 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A2 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A3 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A4 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A5 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_A6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B1 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B2 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B3 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B4 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B5 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_B6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C1 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C2 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C3 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C4 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C5 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_C6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = 1'b0;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D1 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D2 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D3 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D4 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D5 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A1 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A2 = CLBLM_L_X92Y114_SLICE_X145Y114_A5Q;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A4 = CLBLM_L_X92Y113_SLICE_X145Y113_BQ;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A5 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_A6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X155Y134_D6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A1 = CLBLM_L_X98Y133_SLICE_X154Y133_B5Q;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B1 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B2 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B3 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B4 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B5 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_B6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A2 = CLBLL_L_X102Y135_SLICE_X160Y135_CO6;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_A4 = CLBLM_L_X98Y134_SLICE_X154Y134_BO6;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C1 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C2 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C3 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C4 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C5 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_C6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A4 = CLBLL_L_X102Y115_SLICE_X160Y115_CQ;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A5 = CLBLL_L_X102Y115_SLICE_X160Y115_DO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A6 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D1 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D2 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D3 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D4 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D5 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_D6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B1 = CLBLL_L_X102Y115_SLICE_X160Y115_A5Q;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B4 = CLBLL_L_X102Y113_SLICE_X161Y113_DO6;
  assign CLBLM_L_X92Y114_SLICE_X145Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B5 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D1 = CLBLM_L_X98Y134_SLICE_X154Y134_C5Q;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D2 = CLBLM_L_X98Y134_SLICE_X154Y134_AQ;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A1 = CLBLM_L_X92Y114_SLICE_X144Y114_B5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A2 = CLBLM_L_X90Y113_SLICE_X143Y113_A5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A3 = CLBLM_L_X90Y114_SLICE_X143Y114_CO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A4 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_A6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C6 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D3 = CLBLM_R_X97Y132_SLICE_X153Y132_B5Q;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D4 = CLBLM_L_X98Y134_SLICE_X154Y134_A5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B1 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B2 = CLBLM_L_X92Y114_SLICE_X144Y114_BQ;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B3 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B5 = CLBLM_L_X90Y113_SLICE_X143Y113_BQ;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D6 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_B6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D2 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C1 = CLBLM_L_X92Y114_SLICE_X145Y114_AQ;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C2 = CLBLM_R_X93Y119_SLICE_X147Y119_CO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C4 = CLBLM_L_X92Y114_SLICE_X144Y114_A5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C5 = CLBLM_L_X92Y114_SLICE_X144Y114_DO6;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D1 = CLBLM_L_X90Y113_SLICE_X143Y113_BQ;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D2 = CLBLM_R_X93Y114_SLICE_X146Y114_AQ;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D4 = CLBLM_L_X92Y114_SLICE_X144Y114_BQ;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D5 = CLBLM_L_X92Y114_SLICE_X144Y114_B5Q;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_D6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A1 = 1'b1;
  assign CLBLM_L_X92Y114_SLICE_X144Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A2 = CLBLL_L_X102Y114_SLICE_X160Y114_CQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A3 = CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A6 = 1'b1;
  assign LIOB33_X0Y87_IOB_X0Y87_O = 1'b0;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B2 = CLBLL_L_X102Y114_SLICE_X160Y114_CQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B3 = CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B4 = CLBLL_L_X102Y114_SLICE_X160Y114_BQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B6 = CLBLL_L_X102Y114_SLICE_X161Y114_A5Q;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_D1 = CLBLM_R_X93Y125_SLICE_X146Y125_C5Q;
  assign LIOB33_X0Y87_IOB_X0Y87_T = 1'b1;
  assign LIOB33_X0Y87_IOB_X0Y88_T = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y175_IOB_X1Y175_O = 1'b0;
  assign RIOB33_X105Y175_IOB_X1Y176_O = 1'b0;
  assign RIOB33_X105Y175_IOB_X1Y176_T = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_T = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = 1'b0;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A1 = CLBLM_R_X95Y129_SLICE_X151Y129_DQ;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A2 = CLBLM_R_X95Y130_SLICE_X151Y130_C5Q;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A4 = CLBLM_R_X93Y128_SLICE_X147Y128_BQ;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A5 = CLBLM_R_X95Y129_SLICE_X151Y129_B5Q;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_A6 = CLBLM_R_X95Y129_SLICE_X151Y129_BQ;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B2 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B3 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B4 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B5 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_B6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C2 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C3 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C4 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C5 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_C6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = 1'b0;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = 1'b0;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D2 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D3 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D4 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D5 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X151Y128_D6 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = CLBLM_R_X101Y113_SLICE_X159Y113_AO6;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A1 = CLBLM_R_X95Y128_SLICE_X150Y128_B5Q;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A2 = CLBLM_R_X95Y130_SLICE_X150Y130_AQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A3 = CLBLM_R_X95Y128_SLICE_X150Y128_AQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A5 = CLBLM_R_X95Y130_SLICE_X150Y130_CQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_A6 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = 1'b0;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B3 = CLBLM_R_X95Y130_SLICE_X150Y130_CQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B4 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B5 = CLBLM_L_X94Y127_SLICE_X149Y127_BQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = 1'b0;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C1 = CLBLM_R_X95Y130_SLICE_X150Y130_AQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C2 = CLBLM_R_X95Y128_SLICE_X150Y128_AQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C3 = CLBLM_R_X95Y130_SLICE_X150Y130_CQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C4 = CLBLM_R_X93Y128_SLICE_X147Y128_CQ;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C5 = CLBLM_R_X95Y128_SLICE_X150Y128_B5Q;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D1 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D2 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D3 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D4 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D5 = 1'b1;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = 1'b0;
  assign CLBLM_R_X95Y128_SLICE_X150Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A1 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A2 = CLBLM_L_X94Y114_SLICE_X149Y114_AQ;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A3 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A5 = CLBLM_L_X92Y115_SLICE_X145Y115_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_A6 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B1 = CLBLM_L_X92Y115_SLICE_X145Y115_DO6;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B2 = CLBLM_R_X93Y115_SLICE_X147Y115_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B3 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B5 = CLBLM_L_X90Y114_SLICE_X143Y114_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_B6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A1 = CLBLM_R_X101Y116_SLICE_X158Y116_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A2 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A3 = CLBLL_L_X102Y116_SLICE_X160Y116_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A5 = CLBLL_L_X102Y115_SLICE_X160Y115_CO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A6 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_C3 = CLBLM_L_X90Y114_SLICE_X142Y114_DO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B1 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B3 = CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B5 = CLBLL_L_X102Y115_SLICE_X160Y115_BQ;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B6 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D1 = CLBLM_L_X92Y115_SLICE_X145Y115_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C2 = CLBLL_L_X102Y115_SLICE_X160Y115_CQ;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D4 = CLBLM_R_X93Y116_SLICE_X146Y116_CO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C6 = CLBLL_L_X102Y115_SLICE_X161Y115_C5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D5 = CLBLM_L_X94Y116_SLICE_X149Y116_A5Q;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_D6 = CLBLM_L_X90Y114_SLICE_X143Y114_DO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y115_SLICE_X145Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A1 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A2 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_CX = CLBLL_L_X102Y115_SLICE_X161Y115_AO5;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D1 = CLBLL_L_X102Y114_SLICE_X160Y114_C5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D2 = CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D5 = CLBLL_L_X102Y115_SLICE_X160Y115_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_A5 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B4 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B1 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B2 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B5 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_B6 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C1 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C2 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C3 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C4 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C5 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_C6 = 1'b1;
  assign LIOB33_X0Y89_IOB_X0Y89_O = 1'b0;
  assign LIOB33_X0Y89_IOB_X0Y90_T = 1'b1;
  assign LIOB33_X0Y89_IOB_X0Y89_T = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D1 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D2 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A4 = CLBLL_L_X102Y116_SLICE_X161Y116_DO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A5 = CLBLL_L_X102Y116_SLICE_X161Y116_CQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A6 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D4 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D5 = 1'b1;
  assign CLBLM_L_X92Y115_SLICE_X144Y115_D6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B1 = CLBLL_L_X102Y116_SLICE_X160Y116_CQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B5 = CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B6 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y178_O = 1'b0;
  assign RIOB33_X105Y177_IOB_X1Y177_O = 1'b0;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C1 = CLBLL_L_X102Y114_SLICE_X160Y114_C5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C2 = CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C4 = CLBLM_R_X101Y117_SLICE_X158Y117_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C5 = CLBLL_L_X102Y116_SLICE_X161Y116_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y177_IOB_X1Y178_T = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y177_T = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D2 = CLBLL_L_X102Y116_SLICE_X160Y116_CQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D4 = CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D5 = CLBLL_L_X102Y115_SLICE_X161Y115_B5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D6 = CLBLL_L_X102Y116_SLICE_X161Y116_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_X0Y89_IOB_X0Y90_O = 1'b0;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A1 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A3 = CLBLM_R_X95Y129_SLICE_X151Y129_A5Q;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A4 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A5 = CLBLM_R_X95Y126_SLICE_X151Y126_AQ;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_A6 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B1 = CLBLM_L_X98Y129_SLICE_X155Y129_DO6;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B3 = CLBLM_R_X95Y129_SLICE_X151Y129_AQ;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_B6 = CLBLM_R_X95Y129_SLICE_X151Y129_CO6;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_BX = CLBLM_R_X95Y129_SLICE_X151Y129_CO5;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C1 = CLBLM_R_X95Y130_SLICE_X151Y130_C5Q;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C3 = CLBLM_R_X95Y129_SLICE_X151Y129_BQ;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C4 = CLBLM_R_X95Y129_SLICE_X151Y129_DQ;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C5 = CLBLM_R_X95Y129_SLICE_X151Y129_B5Q;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_C6 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D2 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D3 = CLBLM_R_X95Y129_SLICE_X151Y129_BQ;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D4 = CLBLM_R_X95Y129_SLICE_X150Y129_CQ;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D5 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_D6 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X151Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A4 = CLBLM_R_X95Y129_SLICE_X150Y129_BO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A5 = CLBLM_R_X95Y129_SLICE_X151Y129_A5Q;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_A6 = CLBLM_L_X98Y129_SLICE_X154Y129_CO6;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_AX = CLBLM_R_X95Y129_SLICE_X150Y129_BO5;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B1 = CLBLM_R_X95Y129_SLICE_X150Y129_CQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B2 = CLBLM_R_X95Y129_SLICE_X151Y129_D5Q;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B3 = CLBLM_R_X95Y129_SLICE_X150Y129_AQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B5 = CLBLM_R_X95Y129_SLICE_X150Y129_A5Q;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_B6 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C2 = CLBLM_R_X95Y129_SLICE_X150Y129_AQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C3 = CLBLM_L_X94Y129_SLICE_X148Y129_BQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C4 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C5 = 1'b1;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_C6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = 1'b0;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D2 = CLBLM_R_X95Y129_SLICE_X150Y129_AQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D3 = CLBLM_R_X95Y129_SLICE_X151Y129_D5Q;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D4 = CLBLM_R_X95Y129_SLICE_X150Y129_A5Q;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D5 = CLBLM_R_X95Y129_SLICE_X150Y129_CQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_D6 = CLBLM_R_X93Y128_SLICE_X147Y128_AQ;
  assign CLBLM_R_X95Y129_SLICE_X150Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A3 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A1 = CLBLM_L_X92Y116_SLICE_X145Y116_B5Q;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A2 = CLBLM_R_X89Y115_SLICE_X141Y115_CQ;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A3 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A5 = CLBLL_L_X100Y116_SLICE_X157Y116_CO6;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_A6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B1 = CLBLM_L_X90Y116_SLICE_X142Y116_CQ;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B3 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B4 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A3 = CLBLL_L_X102Y116_SLICE_X160Y116_AQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A4 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A4 = CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A5 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_A6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B5 = CLBLM_L_X92Y116_SLICE_X145Y116_BQ;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_B6 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_AX = CLBLM_R_X101Y116_SLICE_X159Y116_AO5;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B1 = CLBLM_R_X101Y116_SLICE_X158Y116_A5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B2 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B3 = CLBLL_L_X102Y116_SLICE_X161Y116_CO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B5 = CLBLL_L_X102Y116_SLICE_X160Y116_C5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_B6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_C5 = CLBLM_L_X92Y116_SLICE_X145Y116_DO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C1 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C2 = CLBLL_L_X100Y117_SLICE_X156Y117_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C3 = CLBLL_L_X100Y117_SLICE_X157Y117_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C5 = CLBLL_L_X102Y116_SLICE_X160Y116_DO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_C6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D1 = CLBLM_L_X90Y116_SLICE_X142Y116_AQ;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D2 = CLBLM_L_X90Y116_SLICE_X142Y116_CQ;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D4 = CLBLM_L_X92Y116_SLICE_X145Y116_BQ;
  assign CLBLM_L_X92Y116_SLICE_X145Y116_D5 = CLBLM_L_X92Y116_SLICE_X145Y116_B5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A1 = CLBLM_L_X90Y118_SLICE_X142Y118_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D2 = CLBLL_L_X102Y116_SLICE_X160Y116_AQ;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D3 = CLBLM_R_X101Y117_SLICE_X158Y117_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D4 = CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_D6 = CLBLL_L_X100Y117_SLICE_X156Y117_DO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A3 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A2 = CLBLM_L_X92Y119_SLICE_X144Y119_CQ;
  assign CLBLL_L_X102Y116_SLICE_X160Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B3 = CLBLM_L_X92Y116_SLICE_X144Y116_AQ;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B4 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B5 = CLBLM_L_X92Y116_SLICE_X144Y116_BQ;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B1 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_A6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C1 = CLBLM_R_X93Y120_SLICE_X146Y120_DO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C2 = CLBLM_L_X90Y116_SLICE_X143Y116_AQ;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C3 = CLBLM_L_X90Y116_SLICE_X143Y116_C5Q;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C5 = CLBLM_L_X92Y116_SLICE_X144Y116_DO6;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = 1'b0;
  assign RIOB33_X105Y179_IOB_X1Y180_O = 1'b0;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A2 = CLBLL_L_X102Y115_SLICE_X161Y115_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A3 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A4 = CLBLL_L_X102Y116_SLICE_X160Y116_BQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A5 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_A6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_D2 = CLBLM_L_X92Y116_SLICE_X144Y116_AQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B2 = CLBLL_L_X102Y116_SLICE_X161Y116_BQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B3 = CLBLL_L_X102Y116_SLICE_X161Y116_AQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B4 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B5 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_B6 = 1'b1;
  assign CLBLM_L_X92Y116_SLICE_X144Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C2 = CLBLL_L_X102Y116_SLICE_X161Y116_CQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C3 = CLBLL_L_X100Y116_SLICE_X156Y116_DO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C4 = CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C5 = CLBLL_L_X102Y116_SLICE_X161Y116_DO6;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A2 = CLBLM_R_X93Y123_SLICE_X146Y123_AQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_CX = CLBLL_L_X102Y116_SLICE_X160Y116_AO5;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D2 = CLBLL_L_X102Y116_SLICE_X161Y116_AQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D3 = CLBLL_L_X102Y116_SLICE_X161Y116_BQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D4 = 1'b1;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D5 = CLBLL_L_X102Y116_SLICE_X161Y116_B5Q;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_D6 = CLBLL_L_X102Y116_SLICE_X160Y116_BQ;
  assign CLBLL_L_X102Y116_SLICE_X161Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B1 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B2 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B3 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A1 = CLBLM_R_X95Y131_SLICE_X150Y131_B5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A2 = CLBLM_L_X98Y131_SLICE_X154Y131_DO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A4 = CLBLM_R_X95Y130_SLICE_X151Y130_BO6;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_AX = CLBLM_R_X95Y130_SLICE_X151Y130_BO5;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B1 = CLBLM_R_X95Y130_SLICE_X151Y130_AQ;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B2 = CLBLM_R_X95Y130_SLICE_X151Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B3 = CLBLM_R_X95Y130_SLICE_X151Y130_CQ;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B4 = CLBLM_R_X95Y131_SLICE_X151Y131_D5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_B6 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C5 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C2 = CLBLM_R_X95Y129_SLICE_X151Y129_DQ;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C3 = CLBLM_R_X95Y130_SLICE_X151Y130_AQ;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C4 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C5 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_C6 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D1 = CLBLM_R_X95Y130_SLICE_X151Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D2 = CLBLM_R_X95Y130_SLICE_X151Y130_CQ;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D4 = CLBLM_R_X93Y128_SLICE_X147Y128_B5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D5 = CLBLM_R_X95Y130_SLICE_X151Y130_AQ;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_D6 = CLBLM_R_X95Y131_SLICE_X151Y131_D5Q;
  assign CLBLM_R_X95Y130_SLICE_X151Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A1 = CLBLM_L_X98Y130_SLICE_X154Y130_DO6;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A4 = CLBLM_L_X94Y130_SLICE_X149Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A5 = CLBLM_R_X95Y128_SLICE_X150Y128_AO6;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_AX = CLBLM_R_X95Y130_SLICE_X150Y130_BO5;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B1 = CLBLM_R_X95Y131_SLICE_X150Y131_CQ;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B2 = CLBLM_R_X95Y130_SLICE_X150Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B4 = CLBLM_R_X95Y132_SLICE_X150Y132_BQ;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B5 = CLBLM_R_X95Y130_SLICE_X150Y130_C5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_B6 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C2 = CLBLM_R_X95Y130_SLICE_X150Y130_AQ;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C3 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C4 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C5 = CLBLM_R_X95Y132_SLICE_X150Y132_BQ;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_C6 = 1'b1;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D1 = CLBLM_R_X95Y130_SLICE_X150Y130_C5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D2 = CLBLM_R_X95Y131_SLICE_X150Y131_CQ;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D3 = CLBLM_R_X93Y131_SLICE_X147Y131_B5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D4 = CLBLM_R_X95Y130_SLICE_X150Y130_A5Q;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_D6 = CLBLM_R_X95Y132_SLICE_X150Y132_BQ;
  assign CLBLM_R_X95Y130_SLICE_X150Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X98Y115_SLICE_X154Y115_B5 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = 1'b0;
  assign LIOB33_X0Y93_IOB_X0Y94_O = 1'b0;
  assign LIOB33_X0Y93_IOB_X0Y93_O = 1'b0;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A1 = CLBLL_L_X102Y117_SLICE_X160Y117_DO6;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A3 = CLBLL_L_X102Y117_SLICE_X161Y117_C5Q;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_A6 = CLBLL_L_X100Y119_SLICE_X156Y119_CO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOB33_X0Y93_IOB_X0Y93_T = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B1 = CLBLL_L_X102Y117_SLICE_X160Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B3 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B4 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B5 = CLBLM_R_X101Y117_SLICE_X159Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_B6 = 1'b1;
  assign LIOB33_X0Y93_IOB_X0Y94_T = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = 1'b0;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C1 = CLBLM_R_X101Y117_SLICE_X159Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C2 = CLBLL_L_X102Y117_SLICE_X160Y117_AQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C4 = CLBLL_L_X102Y117_SLICE_X160Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C5 = CLBLL_L_X102Y117_SLICE_X160Y117_B5Q;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_C6 = CLBLL_L_X102Y117_SLICE_X161Y117_C5Q;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_D1 = 1'b0;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D1 = CLBLM_R_X101Y117_SLICE_X159Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D2 = CLBLL_L_X102Y117_SLICE_X160Y117_AQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D3 = CLBLL_L_X102Y117_SLICE_X160Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D5 = CLBLL_L_X102Y117_SLICE_X160Y117_B5Q;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_D6 = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y181_O = 1'b0;
  assign CLBLL_L_X102Y117_SLICE_X160Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLM_R_X103Y121_SLICE_X162Y121_CO6;
  assign RIOB33_X105Y181_IOB_X1Y182_T = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y181_T = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_D1 = 1'b0;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = 1'b0;
  assign LIOI3_X0Y67_OLOGIC_X0Y67_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = CLBLM_R_X101Y113_SLICE_X159Y113_BO6;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A1 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A2 = CLBLL_L_X102Y117_SLICE_X161Y117_BQ;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A3 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A5 = CLBLL_L_X102Y117_SLICE_X161Y117_A5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = 1'b0;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B1 = CLBLL_L_X102Y117_SLICE_X161Y117_B5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B3 = CLBLL_L_X102Y117_SLICE_X161Y117_CQ;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B4 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B5 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = 1'b0;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C2 = CLBLL_L_X102Y122_SLICE_X160Y122_BQ;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C3 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C4 = CLBLL_L_X102Y117_SLICE_X161Y117_C5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C5 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = 1'b0;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D2 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D3 = CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D4 = CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D5 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLL_L_X102Y117_SLICE_X161Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A1 = CLBLM_R_X95Y131_SLICE_X150Y131_BQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A2 = CLBLM_R_X97Y131_SLICE_X153Y131_DO6;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A4 = CLBLM_R_X95Y131_SLICE_X151Y131_BO6;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_AX = CLBLM_R_X95Y131_SLICE_X151Y131_BO5;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B1 = CLBLM_R_X95Y131_SLICE_X151Y131_AQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B2 = CLBLM_R_X95Y131_SLICE_X151Y131_A5Q;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B4 = CLBLM_R_X95Y131_SLICE_X151Y131_DQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B5 = CLBLM_R_X95Y131_SLICE_X151Y131_C5Q;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_B6 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C2 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C3 = CLBLM_R_X95Y131_SLICE_X151Y131_DQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C4 = CLBLM_R_X97Y131_SLICE_X153Y131_AQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C5 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_C6 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D2 = CLBLM_R_X95Y130_SLICE_X151Y130_CQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D3 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D4 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D5 = CLBLM_R_X95Y131_SLICE_X151Y131_AQ;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_D6 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X151Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A1 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A2 = CLBLM_R_X95Y131_SLICE_X150Y131_BQ;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A4 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A5 = CLBLM_R_X95Y131_SLICE_X150Y131_A5Q;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_A6 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B1 = CLBLM_R_X95Y131_SLICE_X150Y131_B5Q;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B2 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B4 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B5 = CLBLM_R_X95Y129_SLICE_X151Y129_AQ;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_B6 = 1'b1;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C2 = CLBLM_R_X95Y130_SLICE_X150Y130_BO6;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C4 = CLBLM_R_X95Y132_SLICE_X151Y132_AQ;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C5 = CLBLM_R_X97Y133_SLICE_X152Y133_DO6;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y95_IOB_X0Y96_O = 1'b0;
  assign LIOB33_X0Y95_IOB_X0Y95_O = 1'b0;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D1 = CLBLM_R_X93Y129_SLICE_X147Y129_AQ;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D2 = CLBLM_R_X95Y131_SLICE_X151Y131_A5Q;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D3 = CLBLM_R_X95Y131_SLICE_X151Y131_AQ;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D5 = CLBLM_R_X95Y131_SLICE_X151Y131_DQ;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_D6 = CLBLM_R_X95Y131_SLICE_X151Y131_C5Q;
  assign CLBLM_R_X95Y131_SLICE_X150Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y95_IOB_X0Y95_T = 1'b1;
  assign LIOB33_X0Y95_IOB_X0Y96_T = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A2 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A3 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_A4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A2 = CLBLM_R_X101Y118_SLICE_X159Y118_CQ;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A5 = CLBLM_R_X101Y118_SLICE_X159Y118_DO6;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_A6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_B6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B3 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B4 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_B5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_C6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C2 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C3 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C4 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C5 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_C6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X160Y118_D6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D3 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X145Y118_D6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A2 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A3 = CLBLM_R_X89Y115_SLICE_X141Y115_BQ;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A5 = CLBLM_L_X92Y119_SLICE_X144Y119_AQ;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOB33_X105Y97_IOB_X1Y98_O = CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  assign RIOB33_X105Y97_IOB_X1Y97_O = CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B2 = CLBLM_R_X89Y118_SLICE_X141Y118_A5Q;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B3 = CLBLM_R_X89Y115_SLICE_X141Y115_BQ;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B4 = CLBLM_R_X89Y118_SLICE_X141Y118_AQ;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B5 = CLBLM_R_X97Y119_SLICE_X152Y119_CQ;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_B6 = CLBLM_L_X92Y118_SLICE_X144Y118_A5Q;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C2 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C3 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_A6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C5 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_C6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_B6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D1 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_D2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_C6 = 1'b1;
  assign CLBLM_L_X92Y118_SLICE_X144Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D1 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D2 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D3 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D4 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D5 = 1'b1;
  assign CLBLL_L_X102Y118_SLICE_X161Y118_D6 = 1'b1;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C4 = CLBLM_R_X95Y125_SLICE_X151Y125_A5Q;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y124_SLICE_X150Y124_C6 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A1 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A2 = CLBLM_R_X95Y132_SLICE_X151Y132_A5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A4 = CLBLM_R_X97Y132_SLICE_X152Y132_AQ;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A5 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_A6 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B1 = CLBLM_L_X98Y132_SLICE_X154Y132_DO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B3 = CLBLM_R_X95Y132_SLICE_X150Y132_AO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_B6 = CLBLM_R_X95Y132_SLICE_X151Y132_A5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_BX = CLBLM_R_X95Y132_SLICE_X151Y132_DO5;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B1 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C4 = CLBLM_L_X98Y134_SLICE_X154Y134_DO6;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B2 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C5 = CLBLM_R_X95Y132_SLICE_X151Y132_DO6;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_C6 = CLBLM_R_X97Y132_SLICE_X152Y132_AQ;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B4 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D2 = CLBLM_R_X95Y132_SLICE_X151Y132_CQ;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D3 = CLBLM_R_X97Y132_SLICE_X152Y132_DQ;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D4 = CLBLM_R_X95Y132_SLICE_X150Y132_C5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D5 = CLBLM_R_X95Y132_SLICE_X151Y132_B5Q;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_D6 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X151Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A1 = CLBLM_R_X95Y132_SLICE_X150Y132_CQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A2 = CLBLM_R_X95Y132_SLICE_X150Y132_B5Q;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A4 = CLBLM_R_X95Y132_SLICE_X151Y132_BQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A5 = CLBLM_R_X95Y132_SLICE_X150Y132_AQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_A6 = 1'b1;
  assign LIOB33_X0Y97_IOB_X0Y97_O = 1'b0;
  assign LIOB33_X0Y97_IOB_X0Y98_O = 1'b0;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = 1'b0;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B1 = CLBLM_R_X95Y132_SLICE_X150Y132_CQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B2 = CLBLM_R_X95Y131_SLICE_X150Y131_CQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B4 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B5 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_B6 = 1'b1;
  assign LIOB33_X0Y97_IOB_X0Y97_T = 1'b1;
  assign LIOB33_X0Y97_IOB_X0Y98_T = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C2 = CLBLM_R_X97Y132_SLICE_X152Y132_DQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C3 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C4 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C5 = CLBLM_R_X95Y132_SLICE_X151Y132_BQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_C6 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D1 = CLBLM_R_X93Y131_SLICE_X147Y131_BQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D2 = CLBLM_R_X95Y132_SLICE_X150Y132_CQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D3 = CLBLM_R_X95Y132_SLICE_X150Y132_AQ;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C5 = 1'b1;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D5 = CLBLM_R_X95Y132_SLICE_X150Y132_B5Q;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_D6 = CLBLM_R_X95Y132_SLICE_X151Y132_BQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C5 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y185_O = 1'b0;
  assign CLBLM_R_X95Y132_SLICE_X150Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y185_IOB_X1Y186_O = 1'b0;
  assign RIOB33_X105Y185_IOB_X1Y186_T = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y185_T = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A1 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A2 = CLBLM_L_X92Y119_SLICE_X145Y119_A5Q;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A2 = CLBLL_L_X102Y119_SLICE_X161Y119_B5Q;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A3 = CLBLM_L_X92Y115_SLICE_X145Y115_AQ;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A6 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A5 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_A6 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A3 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A4 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_A5 = CLBLL_L_X102Y120_SLICE_X160Y120_AQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B1 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B3 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B4 = CLBLM_L_X90Y119_SLICE_X143Y119_BQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B5 = CLBLM_L_X92Y119_SLICE_X145Y119_BQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_B6 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_B2 = CLBLL_L_X102Y119_SLICE_X160Y119_BQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C1 = CLBLM_L_X92Y118_SLICE_X144Y118_AQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C2 = CLBLM_L_X92Y120_SLICE_X145Y120_C5Q;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C4 = CLBLM_R_X97Y120_SLICE_X153Y120_C5Q;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C5 = CLBLM_L_X92Y119_SLICE_X144Y119_AQ;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C1 = CLBLL_L_X102Y120_SLICE_X160Y120_AQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_C6 = CLBLM_L_X92Y119_SLICE_X144Y119_A5Q;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C2 = CLBLM_R_X103Y120_SLICE_X162Y120_CQ;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C3 = CLBLL_L_X102Y119_SLICE_X160Y119_AQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C4 = CLBLL_L_X102Y119_SLICE_X160Y119_BQ;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C5 = CLBLL_L_X102Y119_SLICE_X160Y119_B5Q;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D1 = CLBLM_R_X93Y124_SLICE_X147Y124_AQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D4 = CLBLM_L_X92Y119_SLICE_X145Y119_BQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D3 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D1 = CLBLL_L_X102Y120_SLICE_X160Y120_AQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D5 = CLBLM_L_X92Y119_SLICE_X145Y119_B5Q;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_D6 = CLBLM_L_X90Y119_SLICE_X143Y119_BQ;
  assign CLBLM_L_X92Y119_SLICE_X145Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D3 = CLBLL_L_X102Y119_SLICE_X160Y119_BQ;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D5 = CLBLL_L_X102Y119_SLICE_X160Y119_B5Q;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y119_SLICE_X160Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A3 = CLBLM_L_X92Y119_SLICE_X144Y119_BO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A5 = CLBLM_L_X90Y123_SLICE_X143Y123_DO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_A6 = CLBLM_L_X92Y121_SLICE_X144Y121_A5Q;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_AX = CLBLM_L_X92Y119_SLICE_X144Y119_BO5;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B1 = CLBLM_L_X92Y118_SLICE_X144Y118_AQ;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B3 = CLBLM_L_X92Y119_SLICE_X144Y119_AQ;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B4 = CLBLM_L_X92Y120_SLICE_X145Y120_C5Q;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B5 = CLBLM_L_X92Y119_SLICE_X144Y119_A5Q;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_B6 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = 1'b0;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C1 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A2 = CLBLM_R_X101Y120_SLICE_X158Y120_DO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C2 = CLBLM_L_X92Y116_SLICE_X144Y116_CO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C3 = CLBLM_L_X92Y119_SLICE_X145Y119_B5Q;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C5 = CLBLM_L_X90Y120_SLICE_X143Y120_A5Q;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_C6 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A4 = CLBLL_L_X102Y119_SLICE_X161Y119_DO6;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A5 = CLBLM_R_X103Y120_SLICE_X162Y120_C5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B2 = CLBLL_L_X102Y119_SLICE_X161Y119_BQ;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B3 = CLBLL_L_X102Y119_SLICE_X161Y119_AQ;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B4 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_B5 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D1 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D2 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D3 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D6 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D4 = 1'b1;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_D5 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C1 = CLBLL_L_X102Y119_SLICE_X161Y119_BQ;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C2 = CLBLL_L_X102Y119_SLICE_X160Y119_A5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C3 = CLBLM_R_X103Y120_SLICE_X162Y120_C5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C5 = CLBLL_L_X102Y119_SLICE_X161Y119_B5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_C6 = CLBLL_L_X102Y119_SLICE_X161Y119_AQ;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y119_SLICE_X144Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D1 = CLBLL_L_X102Y119_SLICE_X161Y119_BQ;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D2 = CLBLL_L_X102Y119_SLICE_X160Y119_A5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D3 = 1'b1;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D5 = CLBLL_L_X102Y119_SLICE_X161Y119_B5Q;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_D6 = CLBLL_L_X102Y119_SLICE_X161Y119_AQ;
  assign CLBLL_L_X102Y119_SLICE_X161Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = 1'b0;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_D1 = CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = 1'b0;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_D1 = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B1 = CLBLM_R_X89Y128_SLICE_X140Y128_AQ;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B2 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B2 = CLBLM_R_X89Y128_SLICE_X140Y128_A5Q;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B6 = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y72_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C6 = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = 1'b0;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D6 = 1'b1;
  assign LIOI3_X0Y71_OLOGIC_X0Y71_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A3 = CLBLM_R_X103Y111_SLICE_X162Y111_AQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A5 = CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_AX = CLBLM_R_X103Y112_SLICE_X162Y112_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B4 = CLBLM_R_X101Y111_SLICE_X159Y111_BQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B5 = CLBLM_R_X103Y111_SLICE_X162Y111_BQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C1 = CLBLM_R_X103Y112_SLICE_X162Y112_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C4 = CLBLM_R_X103Y111_SLICE_X162Y111_BQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C5 = CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C6 = CLBLM_R_X101Y111_SLICE_X159Y111_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = 1'b0;
  assign LIOB33_X0Y101_IOB_X0Y102_O = 1'b0;
  assign LIOB33_X0Y101_IOB_X0Y101_O = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D6 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y101_T = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_T = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y187_IOB_X1Y188_O = 1'b0;
  assign RIOB33_X105Y187_IOB_X1Y187_O = 1'b0;
  assign RIOB33_X105Y187_IOB_X1Y188_T = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_T = 1'b1;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A2 = CLBLL_L_X102Y121_SLICE_X160Y121_BO6;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A4 = CLBLM_R_X103Y120_SLICE_X162Y120_CQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_A6 = CLBLL_L_X102Y119_SLICE_X160Y119_DO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A1 = CLBLM_L_X92Y121_SLICE_X145Y121_DO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B2 = CLBLL_L_X102Y120_SLICE_X160Y120_DQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B3 = CLBLM_R_X101Y117_SLICE_X159Y117_CQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B4 = CLBLM_R_X103Y120_SLICE_X163Y120_B5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_AX = CLBLM_L_X92Y120_SLICE_X145Y120_BO5;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B5 = CLBLM_R_X103Y119_SLICE_X163Y119_B5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B1 = CLBLM_L_X92Y120_SLICE_X145Y120_CQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_B6 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_A4 = CLBLM_L_X92Y120_SLICE_X145Y120_BO6;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B4 = CLBLM_L_X94Y121_SLICE_X148Y121_C5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C1 = CLBLL_L_X102Y119_SLICE_X160Y119_A5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C2 = CLBLL_L_X102Y120_SLICE_X160Y120_CQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C4 = CLBLL_L_X102Y120_SLICE_X160Y120_BQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C5 = CLBLL_L_X102Y119_SLICE_X160Y119_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_C6 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_B3 = CLBLM_L_X92Y120_SLICE_X145Y120_AQ;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C3 = CLBLM_L_X92Y118_SLICE_X144Y118_AQ;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C5 = CLBLM_L_X92Y120_SLICE_X145Y120_AQ;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C6 = 1'b1;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_C1 = 1'b1;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D1 = CLBLL_L_X102Y120_SLICE_X160Y120_C5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D2 = CLBLL_L_X102Y121_SLICE_X161Y121_A5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D4 = CLBLL_L_X102Y120_SLICE_X161Y120_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D5 = CLBLL_L_X102Y120_SLICE_X160Y120_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_D6 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D1 = CLBLM_R_X97Y120_SLICE_X153Y120_CQ;
  assign CLBLL_L_X102Y120_SLICE_X160Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D2 = CLBLM_L_X92Y120_SLICE_X145Y120_CQ;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D4 = CLBLM_L_X92Y120_SLICE_X145Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D5 = CLBLM_L_X92Y120_SLICE_X145Y120_AQ;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_D6 = CLBLM_L_X94Y121_SLICE_X148Y121_C5Q;
  assign CLBLM_L_X92Y120_SLICE_X145Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A1 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A2 = CLBLM_L_X92Y120_SLICE_X144Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A3 = CLBLM_L_X90Y120_SLICE_X142Y120_AQ;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A5 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_A6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B1 = CLBLM_R_X93Y120_SLICE_X146Y120_AQ;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B3 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B4 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B5 = CLBLM_L_X92Y120_SLICE_X144Y120_BQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A2 = CLBLM_R_X103Y120_SLICE_X162Y120_A5Q;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A4 = CLBLL_L_X102Y120_SLICE_X161Y120_DO6;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_A6 = CLBLM_L_X98Y121_SLICE_X155Y121_DO6;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_B6 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C4 = CLBLM_L_X92Y120_SLICE_X144Y120_A5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B2 = CLBLL_L_X102Y120_SLICE_X161Y120_BQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B3 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B4 = 1'b1;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B5 = CLBLL_L_X102Y121_SLICE_X161Y121_AQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_B6 = 1'b1;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C1 = CLBLL_L_X102Y121_SLICE_X161Y121_AQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C3 = CLBLM_R_X103Y120_SLICE_X162Y120_A5Q;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C4 = CLBLL_L_X102Y120_SLICE_X161Y120_BQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C5 = CLBLL_L_X102Y120_SLICE_X161Y120_AQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_C6 = CLBLL_L_X102Y120_SLICE_X161Y120_B5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D1 = CLBLM_L_X92Y120_SLICE_X144Y120_BQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D2 = 1'b1;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D3 = CLBLM_R_X93Y120_SLICE_X146Y120_AQ;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D4 = CLBLM_L_X90Y122_SLICE_X143Y122_C5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D5 = CLBLM_L_X92Y120_SLICE_X144Y120_B5Q;
  assign CLBLM_L_X92Y120_SLICE_X144Y120_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D1 = CLBLL_L_X102Y121_SLICE_X161Y121_AQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D3 = CLBLL_L_X102Y120_SLICE_X161Y120_BQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D4 = CLBLL_L_X102Y120_SLICE_X161Y120_AQ;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D5 = CLBLL_L_X102Y120_SLICE_X161Y120_B5Q;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_D6 = 1'b1;
  assign CLBLL_L_X102Y120_SLICE_X161Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A3 = CLBLM_R_X103Y112_SLICE_X163Y112_AQ;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A5 = CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B3 = CLBLM_R_X103Y112_SLICE_X163Y112_AQ;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B4 = CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B5 = CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B6 = CLBLM_R_X103Y112_SLICE_X163Y112_A5Q;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_BX = CLBLM_R_X103Y113_SLICE_X163Y113_BO5;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y103_IOB_X0Y104_O = 1'b0;
  assign LIOB33_X0Y103_IOB_X0Y103_O = 1'b0;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A1 = CLBLM_R_X103Y112_SLICE_X163Y112_BO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A4 = CLBLM_R_X103Y112_SLICE_X163Y112_BQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_T = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B4 = CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B5 = CLBLM_R_X101Y111_SLICE_X159Y111_AQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y103_T = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C1 = CLBLM_R_X103Y112_SLICE_X162Y112_BQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C2 = CLBLM_R_X103Y112_SLICE_X162Y112_CQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y189_IOB_X1Y190_O = 1'b0;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D1 = CLBLM_R_X103Y112_SLICE_X162Y112_BQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D2 = CLBLM_R_X103Y112_SLICE_X162Y112_CQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D3 = CLBLM_R_X101Y111_SLICE_X159Y111_AQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D4 = CLBLM_R_X103Y112_SLICE_X162Y112_C5Q;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y189_O = 1'b0;
  assign CLBLM_L_X90Y121_SLICE_X143Y121_B6 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A1 = CLBLM_L_X90Y116_SLICE_X143Y116_BQ;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A2 = CLBLM_L_X90Y114_SLICE_X142Y114_C5Q;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A3 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A5 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_A6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y189_IOB_X1Y189_T = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_T = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B1 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B3 = CLBLM_R_X89Y114_SLICE_X141Y114_AQ;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B4 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B5 = CLBLM_R_X89Y114_SLICE_X141Y114_BQ;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_B6 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C1 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C3 = CLBLM_R_X89Y114_SLICE_X141Y114_BQ;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C4 = CLBLM_L_X90Y116_SLICE_X143Y116_BQ;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C5 = CLBLM_R_X89Y114_SLICE_X141Y114_B5Q;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_C6 = CLBLM_R_X89Y114_SLICE_X141Y114_AQ;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D1 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D2 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D3 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D4 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D5 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_D6 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X141Y114_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A1 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A2 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A3 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A4 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A5 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_A6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A2 = CLBLM_R_X101Y120_SLICE_X158Y120_CQ;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A3 = CLBLL_L_X102Y121_SLICE_X160Y121_AQ;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B3 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B4 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B5 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_B6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A4 = CLBLL_L_X100Y121_SLICE_X157Y121_BQ;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A5 = CLBLL_L_X100Y121_SLICE_X157Y121_C5Q;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_A6 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C1 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C2 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C3 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A5 = CLBLM_L_X92Y121_SLICE_X144Y121_CQ;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C4 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A6 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C5 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_C6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C1 = CLBLM_R_X103Y125_SLICE_X162Y125_DO6;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A3 = CLBLM_L_X92Y121_SLICE_X145Y121_AQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_B6 = CLBLM_R_X101Y120_SLICE_X158Y120_CQ;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D1 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D2 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D3 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C1 = CLBLM_L_X92Y121_SLICE_X144Y121_DQ;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D4 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D5 = 1'b1;
  assign CLBLM_R_X89Y114_SLICE_X140Y114_D6 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C5 = CLBLM_L_X94Y121_SLICE_X148Y121_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_C6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D1 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D2 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D3 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D4 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D5 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_D6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X160Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D1 = CLBLM_L_X92Y121_SLICE_X144Y121_CQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D3 = CLBLM_L_X92Y121_SLICE_X145Y121_BQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D5 = CLBLM_L_X92Y121_SLICE_X145Y121_B5Q;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D6 = CLBLM_L_X92Y121_SLICE_X144Y121_DQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_D4 = CLBLM_L_X92Y121_SLICE_X145Y121_AQ;
  assign CLBLM_L_X92Y121_SLICE_X145Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A1 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A2 = CLBLM_L_X92Y121_SLICE_X144Y121_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A3 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A5 = CLBLM_R_X93Y121_SLICE_X146Y121_AQ;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_A6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A2 = CLBLL_L_X102Y120_SLICE_X161Y120_AQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A3 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B4 = CLBLM_R_X93Y121_SLICE_X146Y121_AQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A4 = CLBLM_R_X103Y121_SLICE_X162Y121_B5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B5 = CLBLM_R_X93Y121_SLICE_X146Y121_BO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A5 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_A6 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C2 = CLBLM_L_X92Y121_SLICE_X145Y121_AO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C3 = CLBLM_L_X90Y114_SLICE_X142Y114_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C5 = CLBLM_L_X90Y125_SLICE_X142Y125_BO6;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_C6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B2 = CLBLL_L_X102Y121_SLICE_X161Y121_BQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B3 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B4 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B5 = CLBLM_R_X103Y121_SLICE_X163Y121_BQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_B6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C2 = CLBLL_L_X102Y121_SLICE_X161Y121_CQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C3 = CLBLM_R_X101Y121_SLICE_X159Y121_A5Q;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C4 = CLBLM_R_X103Y121_SLICE_X163Y121_B5Q;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C5 = CLBLL_L_X102Y121_SLICE_X161Y121_B5Q;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_C6 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D6 = 1'b1;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D1 = CLBLM_L_X92Y119_SLICE_X144Y119_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D2 = CLBLM_L_X92Y120_SLICE_X145Y120_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D4 = CLBLM_R_X93Y117_SLICE_X146Y117_A5Q;
  assign CLBLM_L_X92Y121_SLICE_X144Y121_D5 = CLBLM_L_X92Y122_SLICE_X145Y122_CQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D2 = CLBLM_R_X103Y121_SLICE_X163Y121_BQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D3 = CLBLL_L_X102Y121_SLICE_X161Y121_BQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D4 = 1'b1;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D5 = CLBLL_L_X102Y121_SLICE_X161Y121_B5Q;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_D6 = CLBLM_R_X103Y122_SLICE_X163Y122_BQ;
  assign CLBLL_L_X102Y121_SLICE_X161Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A2 = CLBLM_L_X94Y126_SLICE_X149Y126_AO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A4 = CLBLM_L_X92Y125_SLICE_X145Y125_BO6;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A5 = CLBLM_R_X93Y127_SLICE_X146Y127_AQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A4 = CLBLL_L_X102Y114_SLICE_X161Y114_BO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A5 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B3 = CLBLM_R_X103Y113_SLICE_X163Y113_AQ;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B1 = CLBLM_L_X92Y125_SLICE_X145Y125_AQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B4 = CLBLM_R_X103Y113_SLICE_X162Y113_CO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y105_O = 1'b0;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B2 = CLBLM_L_X92Y125_SLICE_X145Y125_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_BX = CLBLL_L_X102Y114_SLICE_X160Y114_AO5;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C2 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C4 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_T = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B4 = CLBLM_L_X92Y125_SLICE_X145Y125_CQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y105_IOB_X0Y105_T = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B5 = CLBLM_L_X92Y125_SLICE_X145Y125_C5Q;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_B6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D4 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A1 = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A2 = CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = 1'b0;
  assign RIOB33_X105Y191_IOB_X1Y192_O = 1'b0;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B4 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B5 = CLBLM_R_X103Y113_SLICE_X162Y113_BQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_T = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_T = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C1 = CLBLM_R_X103Y113_SLICE_X162Y113_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C2 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C4 = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C5 = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C6 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = 1'b0;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D2 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D4 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A1 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A3 = CLBLM_R_X89Y115_SLICE_X141Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A4 = CLBLM_L_X90Y115_SLICE_X142Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A5 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_A6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = 1'b0;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B1 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B3 = CLBLM_R_X89Y115_SLICE_X141Y115_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B4 = CLBLM_R_X89Y118_SLICE_X141Y118_AQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B5 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C1 = CLBLL_L_X102Y113_SLICE_X160Y113_AQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_B6 = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_D1 = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C2 = CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C1 = CLBLM_R_X89Y116_SLICE_X141Y116_C5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C3 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C4 = CLBLM_R_X93Y117_SLICE_X146Y117_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C5 = CLBLM_R_X89Y115_SLICE_X141Y115_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_C6 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y125_SLICE_X142Y125_C2 = 1'b1;
  assign LIOI3_X0Y73_OLOGIC_X0Y74_T1 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D1 = CLBLM_L_X90Y115_SLICE_X142Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D2 = CLBLM_R_X89Y115_SLICE_X141Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D3 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D4 = CLBLM_R_X89Y115_SLICE_X141Y115_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D5 = CLBLM_R_X89Y115_SLICE_X141Y115_B5Q;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C6 = CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  assign LIOI3_X0Y73_OLOGIC_X0Y73_D1 = 1'b0;
  assign CLBLM_R_X89Y115_SLICE_X141Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A1 = CLBLM_R_X89Y116_SLICE_X140Y116_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A2 = CLBLM_L_X90Y119_SLICE_X143Y119_CO6;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A4 = CLBLM_R_X89Y115_SLICE_X140Y115_BO6;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A2 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A3 = CLBLL_L_X102Y122_SLICE_X160Y122_AQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_AX = CLBLM_R_X89Y115_SLICE_X140Y115_BO5;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A4 = CLBLM_R_X101Y123_SLICE_X159Y123_BQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B1 = CLBLM_R_X89Y115_SLICE_X140Y115_CQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B2 = CLBLM_R_X89Y115_SLICE_X140Y115_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B3 = CLBLM_R_X89Y115_SLICE_X140Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B5 = CLBLM_R_X89Y115_SLICE_X140Y115_C5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_B6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A5 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_A6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C1 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C2 = CLBLM_R_X89Y115_SLICE_X140Y115_CQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C3 = CLBLM_R_X89Y115_SLICE_X140Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C5 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_C6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B5 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_B6 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A1 = CLBLM_L_X92Y122_SLICE_X145Y122_B5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A3 = CLBLM_L_X92Y122_SLICE_X145Y122_AQ;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_A4 = CLBLM_L_X92Y123_SLICE_X145Y123_BQ;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B4 = CLBLM_R_X93Y122_SLICE_X146Y122_AQ;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B5 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_B6 = 1'b1;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D1 = CLBLM_R_X89Y115_SLICE_X140Y115_C5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D2 = CLBLM_R_X89Y115_SLICE_X140Y115_CQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D3 = CLBLM_R_X89Y115_SLICE_X140Y115_AQ;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D4 = CLBLM_R_X89Y115_SLICE_X140Y115_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_D6 = CLBLM_R_X89Y116_SLICE_X141Y116_C5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D1 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D2 = CLBLL_L_X102Y122_SLICE_X161Y122_A5Q;
  assign CLBLM_R_X89Y115_SLICE_X140Y115_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D3 = CLBLL_L_X102Y122_SLICE_X160Y122_AQ;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D4 = CLBLL_L_X102Y122_SLICE_X160Y122_A5Q;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_D6 = CLBLM_R_X101Y123_SLICE_X159Y123_BQ;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_C6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X160Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D1 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D3 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D4 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D2 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D5 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_D6 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X145Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A1 = CLBLM_L_X92Y122_SLICE_X144Y122_B5Q;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A2 = CLBLM_L_X90Y122_SLICE_X142Y122_BQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A3 = CLBLM_L_X92Y122_SLICE_X144Y122_AQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A5 = CLBLM_L_X92Y122_SLICE_X144Y122_BQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_A6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A2 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A3 = CLBLL_L_X102Y122_SLICE_X160Y122_A5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A4 = CLBLM_R_X103Y123_SLICE_X162Y123_CQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A5 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_A6 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B2 = CLBLM_L_X92Y122_SLICE_X144Y122_BQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B1 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_B5 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B2 = CLBLL_L_X102Y122_SLICE_X161Y122_BQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B3 = CLBLL_L_X102Y122_SLICE_X161Y122_AQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B4 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C1 = CLBLM_L_X90Y124_SLICE_X143Y124_C5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B5 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_B6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C1 = CLBLM_R_X101Y122_SLICE_X159Y122_CO6;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C2 = CLBLL_L_X102Y122_SLICE_X160Y122_C5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C4 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C5 = CLBLL_L_X102Y122_SLICE_X161Y122_B5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_C6 = 1'b1;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C5 = CLBLM_L_X90Y119_SLICE_X143Y119_CQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_C6 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D3 = CLBLM_L_X92Y122_SLICE_X144Y122_AQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D4 = CLBLM_L_X92Y122_SLICE_X145Y122_CQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D1 = CLBLM_L_X92Y122_SLICE_X144Y122_BQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D2 = CLBLM_R_X103Y123_SLICE_X162Y123_CQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D3 = CLBLL_L_X102Y122_SLICE_X161Y122_BQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D4 = CLBLL_L_X102Y122_SLICE_X161Y122_AQ;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D5 = CLBLL_L_X102Y122_SLICE_X161Y122_B5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_D6 = 1'b1;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D5 = CLBLM_L_X92Y122_SLICE_X144Y122_B5Q;
  assign CLBLL_L_X102Y122_SLICE_X161Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_D6 = CLBLM_L_X90Y122_SLICE_X142Y122_BQ;
  assign CLBLM_L_X92Y122_SLICE_X144Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y107_IOB_X0Y108_O = 1'b0;
  assign LIOB33_X0Y107_IOB_X0Y107_O = 1'b0;
  assign LIOB33_X0Y107_IOB_X0Y108_T = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y107_T = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X103Y120_SLICE_X163Y120_CO6;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLL_L_X102Y118_SLICE_X160Y118_AO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A1 = CLBLM_R_X89Y116_SLICE_X141Y116_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A2 = CLBLM_R_X89Y116_SLICE_X141Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A3 = CLBLM_R_X89Y116_SLICE_X140Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A5 = CLBLM_R_X89Y116_SLICE_X140Y116_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_T = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B1 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B3 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B4 = CLBLM_R_X89Y116_SLICE_X140Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B5 = CLBLM_R_X89Y116_SLICE_X141Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_B6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_T = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C1 = CLBLM_L_X90Y116_SLICE_X142Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C2 = CLBLM_R_X89Y116_SLICE_X141Y116_CQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C4 = CLBLM_L_X90Y117_SLICE_X142Y117_A5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C5 = CLBLM_R_X89Y118_SLICE_X141Y118_D5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_C6 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D1 = CLBLM_R_X89Y116_SLICE_X141Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D2 = CLBLM_R_X89Y116_SLICE_X141Y116_CQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D3 = CLBLM_R_X89Y116_SLICE_X140Y116_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D5 = CLBLM_R_X89Y116_SLICE_X141Y116_B5Q;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_D6 = CLBLM_R_X89Y116_SLICE_X140Y116_BQ;
  assign CLBLM_R_X89Y116_SLICE_X141Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A1 = CLBLM_R_X89Y117_SLICE_X140Y117_CQ;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A2 = CLBLM_R_X89Y116_SLICE_X140Y116_A5Q;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A2 = CLBLL_L_X102Y123_SLICE_X160Y123_DO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A4 = CLBLL_L_X102Y122_SLICE_X160Y122_B5Q;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_A6 = CLBLM_L_X98Y122_SLICE_X154Y122_CO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A5 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_A6 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B3 = CLBLM_R_X89Y116_SLICE_X141Y116_AO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_B5 = CLBLM_L_X90Y120_SLICE_X142Y120_DO6;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B2 = CLBLL_L_X102Y123_SLICE_X160Y123_BQ;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B3 = CLBLL_L_X102Y124_SLICE_X160Y124_CQ;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B4 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B5 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_BX = CLBLM_R_X89Y116_SLICE_X141Y116_AO5;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_B6 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C1 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C2 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C3 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C4 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C5 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_C6 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C2 = CLBLL_L_X102Y123_SLICE_X160Y123_AQ;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_C3 = CLBLL_L_X102Y123_SLICE_X160Y123_BQ;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B4 = CLBLM_L_X92Y123_SLICE_X145Y123_AQ;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B5 = CLBLM_L_X92Y122_SLICE_X145Y122_AO6;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_B6 = CLBLM_R_X89Y123_SLICE_X140Y123_DO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D1 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_BX = CLBLM_L_X92Y123_SLICE_X145Y123_DO5;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D2 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D3 = 1'b1;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D4 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D5 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C3 = CLBLM_L_X90Y126_SLICE_X142Y126_DO6;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_D6 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C4 = CLBLM_L_X92Y123_SLICE_X145Y123_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C5 = CLBLM_L_X92Y123_SLICE_X145Y123_DO6;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y116_SLICE_X140Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y123_SLICE_X160Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D2 = CLBLM_L_X92Y123_SLICE_X145Y123_CQ;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D3 = CLBLM_R_X93Y122_SLICE_X146Y122_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D4 = CLBLM_R_X93Y123_SLICE_X146Y123_BQ;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D5 = CLBLM_L_X92Y123_SLICE_X145Y123_B5Q;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_D6 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X145Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A1 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A2 = CLBLM_L_X92Y123_SLICE_X144Y123_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A4 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A5 = CLBLM_L_X92Y121_SLICE_X144Y121_AQ;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_A6 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A2 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A3 = CLBLM_R_X101Y124_SLICE_X159Y124_A5Q;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A4 = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B1 = CLBLM_L_X90Y126_SLICE_X143Y126_DO6;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A5 = CLBLL_L_X102Y125_SLICE_X161Y125_C5Q;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_A6 = 1'b1;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B2 = CLBLM_R_X93Y123_SLICE_X146Y123_AO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B4 = CLBLM_L_X92Y123_SLICE_X144Y123_AQ;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_B6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C2 = CLBLM_R_X93Y123_SLICE_X147Y123_AO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C4 = CLBLM_L_X92Y123_SLICE_X144Y123_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C5 = CLBLM_L_X92Y124_SLICE_X144Y124_DO6;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_C6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C3 = CLBLL_L_X102Y123_SLICE_X161Y123_A5Q;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_C6 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D2 = CLBLM_L_X92Y123_SLICE_X144Y123_DQ;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D3 = CLBLM_L_X92Y123_SLICE_X145Y123_B5Q;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D4 = CLBLM_L_X92Y122_SLICE_X145Y122_AQ;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D5 = CLBLM_L_X92Y124_SLICE_X145Y124_A5Q;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_D6 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D5 = 1'b1;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_D6 = CLBLM_R_X101Y124_SLICE_X159Y124_A5Q;
  assign CLBLL_L_X102Y123_SLICE_X161Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y123_SLICE_X144Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y109_IOB_X0Y110_O = 1'b0;
  assign LIOB33_X0Y109_IOB_X0Y109_O = 1'b0;
  assign LIOB33_X0Y109_IOB_X0Y110_T = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y109_T = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_R_X103Y124_SLICE_X162Y124_CO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLL_L_X102Y120_SLICE_X161Y120_CO6;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C4 = CLBLM_L_X94Y125_SLICE_X149Y125_CQ;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C5 = CLBLM_R_X95Y124_SLICE_X151Y124_C5Q;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_C6 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A1 = CLBLM_R_X89Y120_SLICE_X141Y120_DO6;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A3 = CLBLM_R_X89Y117_SLICE_X140Y117_C5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A5 = CLBLM_R_X89Y117_SLICE_X141Y117_BO6;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_AX = CLBLM_R_X89Y117_SLICE_X141Y117_BO5;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B1 = CLBLM_R_X89Y117_SLICE_X141Y117_CQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B2 = CLBLM_R_X89Y117_SLICE_X141Y117_A5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B3 = CLBLM_R_X89Y117_SLICE_X141Y117_AQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B5 = CLBLM_R_X89Y117_SLICE_X141Y117_C5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_B6 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C2 = CLBLM_R_X89Y117_SLICE_X141Y117_CQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C3 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C4 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C5 = CLBLM_R_X89Y117_SLICE_X141Y117_AQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_C6 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X95Y125_SLICE_X150Y125_D3 = CLBLM_R_X95Y125_SLICE_X150Y125_BQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D1 = CLBLM_R_X89Y117_SLICE_X141Y117_C5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D2 = CLBLM_R_X89Y117_SLICE_X141Y117_CQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D3 = CLBLM_R_X89Y117_SLICE_X141Y117_A5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D4 = CLBLM_R_X89Y118_SLICE_X141Y118_D5Q;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D5 = CLBLM_R_X89Y117_SLICE_X141Y117_AQ;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y117_SLICE_X141Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A2 = CLBLL_L_X102Y124_SLICE_X160Y124_A5Q;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A3 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A4 = CLBLM_R_X103Y120_SLICE_X162Y120_AQ;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A2 = CLBLM_R_X89Y117_SLICE_X140Y117_A5Q;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A3 = CLBLM_R_X89Y118_SLICE_X140Y118_AQ;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A5 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A5 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_A6 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_A1 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B1 = CLBLM_L_X90Y119_SLICE_X142Y119_AO6;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B3 = CLBLM_R_X89Y117_SLICE_X141Y117_DO6;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B5 = CLBLM_R_X89Y118_SLICE_X140Y118_AQ;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B4 = CLBLM_L_X98Y123_SLICE_X154Y123_DO6;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_B6 = CLBLL_L_X102Y124_SLICE_X160Y124_A5Q;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C2 = CLBLM_R_X89Y119_SLICE_X140Y119_BQ;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C3 = CLBLM_R_X89Y117_SLICE_X140Y117_C5Q;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C4 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C5 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_C6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C5 = CLBLM_R_X103Y124_SLICE_X163Y124_B5Q;
  assign CLBLL_L_X102Y124_SLICE_X160Y124_C6 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A1 = CLBLM_R_X93Y123_SLICE_X146Y123_CQ;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A4 = CLBLM_L_X92Y124_SLICE_X145Y124_AQ;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A5 = CLBLM_L_X92Y122_SLICE_X145Y122_C5Q;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_A6 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D1 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D2 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D3 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D4 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D5 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_D6 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B5 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_B6 = 1'b1;
  assign CLBLM_R_X89Y117_SLICE_X140Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C1 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C2 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C3 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C4 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_C6 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D1 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D2 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D3 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D4 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D5 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X145Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A2 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A3 = CLBLM_R_X103Y124_SLICE_X162Y124_B5Q;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A4 = CLBLL_L_X102Y124_SLICE_X160Y124_BQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A1 = CLBLM_L_X90Y130_SLICE_X142Y130_DO6;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A4 = CLBLM_L_X92Y124_SLICE_X144Y124_BO6;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A5 = CLBLM_L_X90Y123_SLICE_X142Y123_AQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_A5 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B3 = CLBLL_L_X102Y124_SLICE_X161Y124_AQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_AX = CLBLM_L_X92Y124_SLICE_X144Y124_BO5;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B4 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B1 = CLBLM_L_X92Y124_SLICE_X144Y124_AQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B2 = CLBLM_L_X92Y124_SLICE_X144Y124_A5Q;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B4 = CLBLM_L_X92Y124_SLICE_X144Y124_CQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B5 = CLBLM_L_X92Y124_SLICE_X144Y124_C5Q;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_B6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_B5 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C4 = CLBLL_L_X102Y124_SLICE_X161Y124_AQ;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C5 = CLBLL_L_X102Y124_SLICE_X161Y124_B5Q;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C2 = CLBLM_L_X92Y124_SLICE_X144Y124_CQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C3 = CLBLM_L_X92Y124_SLICE_X144Y124_AQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C4 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C5 = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_C6 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_C6 = CLBLL_L_X102Y124_SLICE_X160Y124_BQ;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D2 = 1'b1;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D3 = CLBLL_L_X102Y124_SLICE_X161Y124_BQ;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D5 = CLBLL_L_X102Y124_SLICE_X161Y124_B5Q;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_D6 = CLBLL_L_X102Y124_SLICE_X160Y124_BQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D1 = CLBLM_L_X92Y124_SLICE_X144Y124_C5Q;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D2 = CLBLM_L_X92Y124_SLICE_X145Y124_AQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D3 = CLBLM_L_X92Y124_SLICE_X144Y124_AQ;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D4 = CLBLM_L_X92Y124_SLICE_X144Y124_A5Q;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_D6 = CLBLM_L_X92Y124_SLICE_X144Y124_CQ;
  assign CLBLL_L_X102Y124_SLICE_X161Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y111_IOB_X0Y111_T = 1'b1;
  assign CLBLM_L_X92Y124_SLICE_X144Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = 1'b0;
  assign LIOI3_X0Y75_OLOGIC_X0Y75_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X103Y124_SLICE_X163Y124_CO6;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLL_L_X102Y124_SLICE_X161Y124_CO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A2 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A3 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A4 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A5 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B2 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B3 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B4 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B5 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C2 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C3 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C4 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C5 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D2 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D3 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D4 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D5 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A2 = CLBLL_L_X102Y117_SLICE_X161Y117_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A4 = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A5 = CLBLM_R_X97Y118_SLICE_X153Y118_DO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B2 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B3 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B4 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B5 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C2 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C3 = CLBLL_L_X102Y117_SLICE_X161Y117_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C4 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C5 = CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C6 = CLBLL_L_X102Y117_SLICE_X161Y117_D5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D2 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D3 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D5 = CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D6 = CLBLL_L_X102Y117_SLICE_X161Y117_D5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A1 = CLBLM_R_X89Y119_SLICE_X141Y119_DO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A4 = CLBLM_R_X89Y118_SLICE_X141Y118_BO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A5 = CLBLM_R_X89Y119_SLICE_X140Y119_AQ;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_AX = CLBLM_R_X89Y118_SLICE_X141Y118_BO5;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B1 = CLBLM_L_X92Y118_SLICE_X144Y118_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B2 = CLBLM_R_X89Y118_SLICE_X141Y118_AQ;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B4 = CLBLM_R_X89Y115_SLICE_X141Y115_BQ;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B5 = CLBLM_R_X89Y118_SLICE_X141Y118_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_B6 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C2 = CLBLM_R_X93Y117_SLICE_X146Y117_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C3 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C4 = CLBLM_R_X89Y118_SLICE_X141Y118_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C5 = CLBLM_R_X89Y120_SLICE_X140Y120_CQ;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_C6 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D1 = CLBLM_L_X90Y119_SLICE_X143Y119_AQ;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D2 = CLBLM_R_X89Y118_SLICE_X141Y118_CQ;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D3 = CLBLM_R_X89Y118_SLICE_X141Y118_DQ;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A2 = CLBLL_L_X102Y126_SLICE_X161Y126_D5Q;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_A6 = CLBLL_L_X102Y125_SLICE_X160Y125_CO6;
  assign CLBLM_R_X89Y118_SLICE_X141Y118_D4 = CLBLM_R_X89Y118_SLICE_X140Y118_B5Q;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A3 = CLBLM_R_X89Y119_SLICE_X140Y119_AQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A4 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_A6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B2 = CLBLL_L_X102Y125_SLICE_X160Y125_BQ;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B3 = CLBLL_L_X102Y125_SLICE_X160Y125_AQ;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B4 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B5 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B2 = CLBLM_R_X89Y118_SLICE_X140Y118_A5Q;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_B6 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_B6 = CLBLM_R_X89Y118_SLICE_X140Y118_CO6;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C1 = CLBLL_L_X102Y126_SLICE_X161Y126_AQ;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C2 = CLBLL_L_X102Y125_SLICE_X160Y125_AQ;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C3 = CLBLL_L_X102Y125_SLICE_X161Y125_B5Q;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_BX = CLBLM_R_X89Y118_SLICE_X140Y118_CO5;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_C4 = CLBLL_L_X102Y125_SLICE_X160Y125_BQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C2 = CLBLM_R_X89Y118_SLICE_X140Y118_B5Q;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C3 = CLBLM_R_X89Y118_SLICE_X140Y118_DQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C4 = CLBLM_L_X90Y118_SLICE_X142Y118_A5Q;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C5 = CLBLM_R_X89Y118_SLICE_X140Y118_BQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_C6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_AX = CLBLM_L_X92Y125_SLICE_X145Y125_BO5;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D1 = CLBLM_R_X101Y126_SLICE_X159Y126_A5Q;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D2 = CLBLL_L_X102Y125_SLICE_X160Y125_AQ;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D3 = CLBLL_L_X102Y125_SLICE_X161Y125_B5Q;
  assign CLBLL_L_X102Y125_SLICE_X160Y125_D4 = CLBLL_L_X102Y125_SLICE_X160Y125_BQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D2 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D3 = CLBLM_L_X92Y122_SLICE_X145Y122_BQ;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D4 = 1'b1;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D5 = CLBLM_R_X89Y118_SLICE_X140Y118_BQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_D6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C2 = CLBLM_L_X92Y125_SLICE_X145Y125_CQ;
  assign CLBLM_R_X89Y118_SLICE_X140Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C5 = CLBLM_L_X92Y125_SLICE_X145Y125_AQ;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_C6 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D1 = CLBLM_L_X92Y125_SLICE_X145Y125_C5Q;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D2 = CLBLM_L_X92Y125_SLICE_X145Y125_CQ;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D4 = CLBLM_L_X92Y125_SLICE_X145Y125_A5Q;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D5 = CLBLM_L_X92Y125_SLICE_X145Y125_AQ;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_D6 = CLBLM_L_X90Y124_SLICE_X143Y124_CQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A1 = CLBLL_L_X102Y125_SLICE_X161Y125_DO6;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A2 = CLBLL_L_X102Y126_SLICE_X160Y126_AQ;
  assign CLBLM_L_X92Y125_SLICE_X145Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_A3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_A6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B2 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_B3 = CLBLL_L_X102Y125_SLICE_X161Y125_AQ;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_B6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C1 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C2 = CLBLL_L_X102Y125_SLICE_X161Y125_CQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_C6 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D1 = CLBLL_L_X102Y125_SLICE_X161Y125_C5Q;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D2 = CLBLL_L_X102Y125_SLICE_X161Y125_CQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D3 = 1'b1;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D4 = CLBLL_L_X102Y125_SLICE_X161Y125_BQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_D6 = CLBLL_L_X102Y125_SLICE_X161Y125_AQ;
  assign CLBLL_L_X102Y125_SLICE_X161Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D1 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D2 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D3 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D4 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D5 = 1'b1;
  assign CLBLM_L_X92Y125_SLICE_X144Y125_D6 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A2 = CLBLL_R_X87Y118_SLICE_X138Y118_BQ;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A3 = CLBLL_R_X87Y118_SLICE_X138Y118_AQ;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A4 = CLBLL_R_X87Y118_SLICE_X138Y118_B5Q;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A5 = CLBLL_R_X87Y118_SLICE_X139Y118_AQ;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_A6 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B1 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B2 = CLBLL_R_X87Y118_SLICE_X138Y118_BQ;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B3 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B5 = CLBLL_R_X87Y118_SLICE_X139Y118_AQ;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_B6 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C1 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C2 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C3 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C4 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C5 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_C6 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D1 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D2 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D3 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D4 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D5 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_D6 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X138Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A2 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A3 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A4 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A6 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B2 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B3 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B4 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B6 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A1 = CLBLM_R_X89Y121_SLICE_X141Y121_DO6;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A3 = CLBLL_R_X87Y118_SLICE_X138Y118_AO6;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A5 = CLBLM_R_X89Y119_SLICE_X140Y119_BQ;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C2 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C3 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B2 = CLBLM_R_X89Y118_SLICE_X141Y118_DQ;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B3 = CLBLL_R_X87Y118_SLICE_X139Y118_AQ;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B4 = CLBLL_R_X87Y118_SLICE_X138Y118_BQ;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B5 = CLBLL_R_X87Y118_SLICE_X138Y118_AQ;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_B6 = CLBLL_R_X87Y118_SLICE_X138Y118_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D2 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C1 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C2 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C3 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C4 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C5 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_C6 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D3 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D4 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A2 = CLBLM_R_X103Y117_SLICE_X162Y117_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A5 = CLBLL_L_X102Y117_SLICE_X161Y117_BQ;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D1 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D2 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D3 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D4 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D5 = 1'b1;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_D6 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A6 = CLBLM_R_X97Y118_SLICE_X152Y118_DO6;
  assign CLBLL_R_X87Y118_SLICE_X139Y118_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B2 = CLBLM_R_X103Y117_SLICE_X162Y117_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B3 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B4 = CLBLL_L_X102Y117_SLICE_X161Y117_DQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B6 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C1 = CLBLL_L_X102Y117_SLICE_X161Y117_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C2 = CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C4 = CLBLM_R_X103Y117_SLICE_X162Y117_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C5 = CLBLM_R_X103Y117_SLICE_X162Y117_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C6 = CLBLL_L_X102Y117_SLICE_X161Y117_DQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D2 = CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D3 = CLBLM_R_X103Y117_SLICE_X162Y117_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D5 = CLBLM_R_X103Y117_SLICE_X162Y117_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D6 = CLBLL_L_X102Y117_SLICE_X161Y117_DQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A4 = CLBLM_R_X89Y119_SLICE_X141Y119_BO6;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A5 = CLBLM_R_X89Y119_SLICE_X140Y119_B5Q;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_A6 = CLBLM_L_X90Y122_SLICE_X143Y122_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_AX = CLBLM_R_X89Y119_SLICE_X141Y119_BO5;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B1 = CLBLM_R_X89Y119_SLICE_X141Y119_AQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B2 = CLBLM_R_X89Y119_SLICE_X141Y119_A5Q;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B4 = CLBLM_R_X89Y119_SLICE_X141Y119_CQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B5 = CLBLM_R_X89Y119_SLICE_X141Y119_C5Q;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_B6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C2 = CLBLM_R_X89Y119_SLICE_X141Y119_CQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C3 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C4 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C5 = CLBLM_R_X89Y119_SLICE_X141Y119_AQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_C6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A2 = CLBLL_L_X102Y126_SLICE_X160Y126_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A3 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D2 = CLBLM_R_X89Y119_SLICE_X141Y119_CQ;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A4 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A5 = CLBLL_L_X102Y126_SLICE_X161Y126_AQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_A6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X141Y119_D1 = CLBLM_R_X89Y119_SLICE_X141Y119_C5Q;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B1 = CLBLL_L_X102Y126_SLICE_X160Y126_DO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B2 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B3 = CLBLL_L_X102Y123_SLICE_X161Y123_DO6;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B5 = CLBLL_L_X102Y126_SLICE_X160Y126_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A1 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A5 = CLBLM_L_X92Y123_SLICE_X145Y123_AQ;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_A2 = CLBLM_R_X89Y119_SLICE_X140Y119_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C1 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C2 = CLBLL_L_X102Y126_SLICE_X160Y126_CQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C4 = CLBLL_L_X102Y126_SLICE_X160Y126_BQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C5 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_C6 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B4 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B5 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B1 = CLBLM_R_X89Y119_SLICE_X140Y119_B5Q;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_B2 = CLBLM_R_X89Y124_SLICE_X140Y124_AQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D2 = CLBLL_L_X102Y126_SLICE_X160Y126_CQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D3 = CLBLL_L_X102Y126_SLICE_X160Y126_BQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D4 = CLBLL_L_X102Y126_SLICE_X160Y126_C5Q;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D5 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_C5 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_D6 = CLBLL_L_X102Y126_SLICE_X161Y126_C5Q;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A1 = CLBLM_L_X92Y126_SLICE_X145Y126_B5Q;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A2 = CLBLM_L_X92Y126_SLICE_X145Y126_BQ;
  assign CLBLL_L_X102Y126_SLICE_X160Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A4 = CLBLM_R_X93Y127_SLICE_X146Y127_CQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A5 = CLBLM_L_X92Y126_SLICE_X144Y126_AQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_A6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B2 = CLBLM_L_X92Y126_SLICE_X145Y126_BQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B3 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B4 = CLBLM_R_X93Y127_SLICE_X146Y127_CQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B5 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C1 = CLBLM_L_X90Y125_SLICE_X143Y125_BQ;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_B6 = CLBLM_L_X94Y124_SLICE_X149Y124_CO6;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C2 = CLBLM_L_X92Y126_SLICE_X145Y126_CQ;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D1 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D2 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D3 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D4 = 1'b1;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D5 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y119_SLICE_X140Y119_D6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C4 = CLBLM_R_X89Y125_SLICE_X141Y125_A5Q;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C5 = CLBLM_R_X89Y126_SLICE_X141Y126_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A2 = CLBLL_L_X102Y126_SLICE_X161Y126_A5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A3 = CLBLL_L_X102Y127_SLICE_X160Y127_AQ;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A4 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A5 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_A6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D1 = CLBLM_L_X92Y126_SLICE_X144Y126_AQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D2 = CLBLM_L_X92Y126_SLICE_X145Y126_CQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D3 = CLBLM_L_X92Y126_SLICE_X145Y126_BQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D4 = CLBLM_R_X93Y127_SLICE_X146Y127_CQ;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A1 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A2 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A3 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A4 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A5 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_A6 = 1'b1;
  assign CLBLM_L_X94Y124_SLICE_X149Y124_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B3 = CLBLM_R_X103Y126_SLICE_X162Y126_AQ;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B4 = CLBLL_L_X102Y127_SLICE_X161Y127_A5Q;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_AX = CLBLM_L_X92Y126_SLICE_X145Y126_AO5;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_B6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B1 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B2 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B3 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B4 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B5 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_B6 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_C4 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D1 = CLBLL_L_X102Y126_SLICE_X161Y126_DQ;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D2 = CLBLL_L_X102Y125_SLICE_X161Y125_B5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D4 = CLBLM_R_X103Y126_SLICE_X162Y126_B5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D5 = CLBLL_L_X102Y127_SLICE_X161Y127_B5Q;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_D6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C1 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C2 = 1'b1;
  assign CLBLL_L_X102Y126_SLICE_X161Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C3 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C4 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C5 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_C6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D1 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D2 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D3 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D4 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D5 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_D6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X144Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y201_OLOGIC_X0Y202_D1 = 1'b0;
  assign LIOI3_X0Y201_OLOGIC_X0Y202_T1 = 1'b1;
  assign LIOI3_X0Y201_OLOGIC_X0Y201_D1 = 1'b0;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_D1 = 1'b0;
  assign LIOI3_X0Y201_OLOGIC_X0Y201_T1 = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y78_T1 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_B6 = 1'b1;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = 1'b0;
  assign LIOI3_X0Y77_OLOGIC_X0Y77_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A1 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A2 = CLBLM_R_X89Y121_SLICE_X141Y121_CQ;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_C6 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A4 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A5 = CLBLM_L_X90Y120_SLICE_X142Y120_BQ;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_A6 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B1 = CLBLM_R_X89Y124_SLICE_X140Y124_CQ;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B2 = CLBLM_R_X89Y119_SLICE_X141Y119_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B4 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B5 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_B6 = CLBLM_L_X90Y115_SLICE_X142Y115_A5Q;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C2 = CLBLM_R_X89Y120_SLICE_X141Y120_CQ;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C3 = CLBLL_R_X87Y118_SLICE_X138Y118_AQ;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C4 = CLBLM_R_X89Y120_SLICE_X141Y120_BQ;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C5 = CLBLM_R_X89Y117_SLICE_X141Y117_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_C6 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A2 = CLBLL_L_X102Y127_SLICE_X160Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A3 = CLBLL_L_X102Y130_SLICE_X161Y130_AQ;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A4 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A5 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_A6 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D1 = CLBLM_R_X89Y120_SLICE_X141Y120_C5Q;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B2 = CLBLL_L_X102Y127_SLICE_X160Y127_DO6;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B4 = CLBLL_L_X102Y127_SLICE_X161Y127_BQ;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D4 = CLBLM_R_X89Y120_SLICE_X141Y120_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X141Y120_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C1 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C2 = CLBLL_L_X102Y127_SLICE_X160Y127_CQ;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A5 = CLBLM_R_X89Y119_SLICE_X140Y119_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C4 = CLBLL_L_X102Y129_SLICE_X160Y129_CQ;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C5 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_AX = CLBLM_R_X89Y120_SLICE_X140Y120_BO5;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_C6 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B1 = CLBLM_R_X89Y118_SLICE_X140Y118_D5Q;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B2 = CLBLM_L_X92Y122_SLICE_X145Y122_BQ;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B4 = CLBLM_R_X89Y120_SLICE_X140Y120_AQ;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B5 = CLBLM_R_X89Y120_SLICE_X140Y120_A5Q;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_B6 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D1 = CLBLL_L_X102Y127_SLICE_X160Y127_C5Q;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D2 = CLBLL_L_X102Y129_SLICE_X160Y129_CQ;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D3 = CLBLL_L_X102Y127_SLICE_X160Y127_BQ;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D4 = CLBLL_L_X102Y127_SLICE_X160Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_D6 = CLBLL_L_X102Y127_SLICE_X160Y127_CQ;
  assign CLBLL_L_X102Y127_SLICE_X160Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D5 = CLBLM_L_X92Y126_SLICE_X145Y126_B5Q;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A4 = CLBLM_L_X92Y127_SLICE_X145Y127_B5Q;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A5 = CLBLM_R_X93Y127_SLICE_X146Y127_BQ;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A6 = 1'b1;
  assign CLBLM_L_X92Y126_SLICE_X145Y126_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B1 = CLBLM_L_X92Y127_SLICE_X145Y127_BQ;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B3 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B4 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B5 = CLBLM_R_X93Y127_SLICE_X146Y127_BQ;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_B6 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D1 = CLBLM_L_X92Y122_SLICE_X145Y122_BQ;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D3 = CLBLM_R_X89Y120_SLICE_X140Y120_AQ;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C1 = CLBLM_R_X93Y127_SLICE_X146Y127_BQ;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D4 = CLBLM_R_X89Y120_SLICE_X140Y120_A5Q;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C2 = CLBLM_L_X90Y125_SLICE_X143Y125_CQ;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_D5 = CLBLM_R_X89Y118_SLICE_X140Y118_D5Q;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C3 = CLBLM_L_X92Y127_SLICE_X145Y127_BQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A2 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A3 = CLBLL_L_X102Y127_SLICE_X161Y127_AQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A4 = CLBLM_R_X103Y127_SLICE_X162Y127_AQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A5 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_A6 = 1'b1;
  assign CLBLM_R_X89Y120_SLICE_X140Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D5 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D6 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B1 = CLBLL_L_X102Y126_SLICE_X161Y126_B5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B2 = CLBLL_L_X102Y127_SLICE_X161Y127_BQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B5 = CLBLL_L_X102Y129_SLICE_X161Y129_AQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_B6 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A1 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C1 = CLBLL_L_X102Y127_SLICE_X160Y127_AQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C2 = CLBLL_L_X102Y126_SLICE_X161Y126_B5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C4 = CLBLL_L_X102Y127_SLICE_X161Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C5 = CLBLL_L_X102Y127_SLICE_X161Y127_AQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_C6 = CLBLM_R_X103Y127_SLICE_X162Y127_AQ;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A2 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A5 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A6 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B1 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B2 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B3 = 1'b1;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D2 = CLBLM_R_X101Y127_SLICE_X159Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D3 = CLBLL_L_X102Y126_SLICE_X161Y126_B5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D4 = CLBLL_L_X102Y127_SLICE_X161Y127_A5Q;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D5 = CLBLL_L_X102Y127_SLICE_X161Y127_AQ;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_D6 = CLBLM_R_X103Y127_SLICE_X162Y127_AQ;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B4 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y127_SLICE_X161Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C1 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B5 = CLBLM_L_X98Y111_SLICE_X155Y111_AQ;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C2 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C3 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C4 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C5 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_B6 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_C6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D1 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D2 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D3 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D4 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D5 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_D6 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C4 = CLBLL_L_X100Y111_SLICE_X156Y111_A5Q;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C5 = CLBLL_L_X100Y111_SLICE_X156Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_C6 = CLBLM_L_X98Y111_SLICE_X155Y111_DO6;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A4 = CLBLM_R_X103Y119_SLICE_X163Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A5 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A6 = CLBLL_L_X100Y119_SLICE_X157Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B2 = CLBLM_R_X103Y119_SLICE_X163Y119_BQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B4 = CLBLM_R_X103Y120_SLICE_X163Y120_BQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C1 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C3 = CLBLM_R_X103Y119_SLICE_X163Y119_BQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C4 = CLBLM_R_X103Y119_SLICE_X163Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C5 = CLBLM_R_X103Y119_SLICE_X163Y119_B5Q;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C6 = CLBLM_R_X103Y120_SLICE_X163Y120_BQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X90Y128_SLICE_X143Y128_D6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D1 = 1'b1;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D3 = CLBLM_R_X103Y119_SLICE_X163Y119_BQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D4 = CLBLM_R_X103Y119_SLICE_X163Y119_AQ;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D5 = CLBLM_R_X103Y119_SLICE_X163Y119_B5Q;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D6 = CLBLM_R_X103Y120_SLICE_X163Y120_BQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y111_SLICE_X156Y111_D4 = CLBLL_L_X100Y111_SLICE_X156Y111_BQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_AX = CLBLL_L_X102Y118_SLICE_X160Y118_AO5;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D6 = 1'b1;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A5 = CLBLM_L_X90Y128_SLICE_X143Y128_CQ;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A1 = CLBLM_R_X93Y125_SLICE_X146Y125_DO6;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A3 = CLBLM_R_X89Y122_SLICE_X141Y122_AQ;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A4 = CLBLM_R_X89Y121_SLICE_X141Y121_BO6;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X90Y128_SLICE_X142Y128_A6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_AX = CLBLM_R_X89Y121_SLICE_X141Y121_BO5;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B1 = CLBLM_R_X89Y121_SLICE_X141Y121_AQ;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B2 = CLBLM_R_X89Y121_SLICE_X141Y121_A5Q;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B4 = CLBLM_R_X89Y120_SLICE_X141Y120_A5Q;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B5 = CLBLM_R_X89Y121_SLICE_X141Y121_CQ;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_B6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = 1'b0;
  assign LIOB33_X0Y119_IOB_X0Y119_O = 1'b0;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C2 = CLBLM_R_X89Y122_SLICE_X141Y122_DQ;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C3 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A1 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A2 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A3 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A4 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_A6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C4 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C5 = CLBLM_R_X89Y121_SLICE_X141Y121_AQ;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_C6 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B1 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B2 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B3 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B4 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_B6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D1 = CLBLM_R_X89Y121_SLICE_X141Y121_C5Q;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C1 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X141Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C2 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C3 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C4 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_C6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A1 = CLBLM_R_X89Y124_SLICE_X140Y124_DO6;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A2 = CLBLM_R_X89Y124_SLICE_X140Y124_AQ;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A4 = CLBLM_R_X89Y121_SLICE_X140Y121_BO6;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_AX = CLBLM_R_X89Y121_SLICE_X140Y121_BO5;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D1 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D2 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D3 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D4 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X160Y128_D6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B1 = CLBLM_R_X89Y121_SLICE_X140Y121_AQ;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B2 = CLBLM_R_X89Y121_SLICE_X140Y121_A5Q;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_B5 = CLBLM_R_X89Y121_SLICE_X140Y121_C5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A2 = CLBLM_L_X94Y129_SLICE_X148Y129_CO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A3 = CLBLM_L_X92Y128_SLICE_X145Y128_BO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A5 = CLBLM_R_X93Y129_SLICE_X146Y129_AQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_AX = CLBLM_L_X92Y128_SLICE_X145Y128_BO5;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_C2 = CLBLM_R_X89Y121_SLICE_X140Y121_CQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B1 = CLBLM_L_X92Y128_SLICE_X145Y128_AQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B2 = CLBLM_L_X92Y128_SLICE_X145Y128_C5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B3 = CLBLM_L_X92Y128_SLICE_X145Y128_A5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B4 = CLBLM_L_X92Y128_SLICE_X145Y128_CQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_B6 = 1'b1;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D1 = CLBLM_R_X89Y121_SLICE_X140Y121_C5Q;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D2 = CLBLM_R_X89Y121_SLICE_X140Y121_CQ;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D3 = CLBLM_R_X89Y121_SLICE_X140Y121_AQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y121_SLICE_X140Y121_D4 = CLBLM_R_X89Y121_SLICE_X140Y121_A5Q;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A2 = CLBLL_L_X102Y129_SLICE_X161Y129_AQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A3 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_A6 = CLBLL_L_X102Y128_SLICE_X161Y128_CO6;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C2 = CLBLM_L_X92Y128_SLICE_X145Y128_CQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C3 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C5 = CLBLM_L_X92Y128_SLICE_X145Y128_AQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B2 = CLBLL_L_X102Y128_SLICE_X161Y128_BQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B3 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B4 = CLBLL_L_X102Y126_SLICE_X161Y126_CQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_B6 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D1 = CLBLM_L_X92Y128_SLICE_X145Y128_C5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D2 = CLBLM_L_X90Y125_SLICE_X143Y125_B5Q;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C1 = CLBLL_L_X102Y128_SLICE_X161Y128_BQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C2 = CLBLL_L_X102Y126_SLICE_X161Y126_CQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C4 = CLBLL_L_X102Y128_SLICE_X161Y128_AQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C5 = CLBLL_L_X102Y128_SLICE_X161Y128_B5Q;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_C6 = CLBLL_L_X102Y130_SLICE_X161Y130_AQ;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A1 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A2 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A3 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A4 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D1 = CLBLL_L_X102Y128_SLICE_X161Y128_BQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D2 = CLBLL_L_X102Y126_SLICE_X161Y126_CQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D4 = CLBLL_L_X102Y128_SLICE_X161Y128_AQ;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B5 = 1'b1;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D6 = CLBLL_L_X100Y129_SLICE_X156Y129_AQ;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_D5 = CLBLL_L_X102Y128_SLICE_X161Y128_B5Q;
  assign CLBLL_L_X102Y128_SLICE_X161Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B2 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B3 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B4 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B6 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C1 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C2 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C3 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C4 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C5 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_C6 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D1 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D2 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D3 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D4 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D5 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_D6 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A1 = CLBLM_R_X103Y120_SLICE_X163Y120_DO6;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A2 = CLBLL_L_X100Y120_SLICE_X157Y120_CO6;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A4 = CLBLM_R_X103Y120_SLICE_X162Y120_BQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B2 = CLBLM_R_X103Y119_SLICE_X163Y119_AQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B3 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B4 = CLBLM_R_X103Y121_SLICE_X163Y121_A5Q;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B5 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_B6 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C1 = CLBLM_R_X103Y121_SLICE_X163Y121_AQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C3 = CLBLM_R_X103Y121_SLICE_X163Y121_A5Q;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C4 = CLBLM_R_X103Y120_SLICE_X163Y120_AQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C5 = CLBLM_R_X103Y120_SLICE_X163Y120_B5Q;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_C6 = CLBLM_R_X103Y120_SLICE_X162Y120_BQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D1 = CLBLM_R_X103Y121_SLICE_X163Y121_AQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D3 = CLBLM_R_X103Y121_SLICE_X163Y121_A5Q;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D4 = CLBLM_R_X103Y120_SLICE_X163Y120_AQ;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D5 = CLBLM_R_X103Y120_SLICE_X163Y120_B5Q;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_D6 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X163Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A2 = CLBLM_R_X103Y120_SLICE_X162Y120_BQ;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A3 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A4 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C2 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A5 = CLBLM_R_X103Y120_SLICE_X162Y120_A5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_A6 = 1'b1;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C3 = CLBLM_R_X95Y126_SLICE_X150Y126_BQ;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B2 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B3 = CLBLM_R_X103Y120_SLICE_X162Y120_CQ;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C4 = CLBLM_R_X95Y126_SLICE_X150Y126_A5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B4 = CLBLM_R_X103Y120_SLICE_X162Y120_B5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B5 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_B6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = 1'b0;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C5 = CLBLM_R_X95Y126_SLICE_X150Y126_B5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C1 = CLBLM_R_X103Y120_SLICE_X162Y120_C5Q;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C2 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X95Y126_SLICE_X150Y126_C6 = CLBLM_R_X97Y126_SLICE_X152Y126_AQ;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C4 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C5 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_C6 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y121_IOB_X0Y122_O = 1'b0;
  assign LIOB33_X0Y121_IOB_X0Y121_O = 1'b0;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D1 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D2 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D3 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D4 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D5 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_T = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A1 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A2 = CLBLM_R_X89Y124_SLICE_X141Y124_AQ;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A4 = CLBLM_R_X89Y122_SLICE_X141Y122_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A5 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y120_SLICE_X162Y120_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y121_IOB_X0Y121_T = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B2 = CLBLM_L_X92Y125_SLICE_X145Y125_DO6;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B3 = CLBLM_R_X89Y122_SLICE_X141Y122_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_B6 = CLBLM_R_X89Y122_SLICE_X141Y122_CO6;
  assign LIOI3_X0Y203_OLOGIC_X0Y204_D1 = 1'b0;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A2 = CLBLL_L_X102Y129_SLICE_X160Y129_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C1 = CLBLM_R_X89Y122_SLICE_X141Y122_BQ;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C3 = CLBLM_R_X89Y122_SLICE_X141Y122_DQ;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C4 = CLBLM_R_X89Y121_SLICE_X141Y121_C5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C5 = CLBLM_R_X89Y122_SLICE_X141Y122_B5Q;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_C6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A3 = CLBLL_L_X100Y128_SLICE_X156Y128_AQ;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A4 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A5 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_A6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B2 = CLBLL_L_X102Y130_SLICE_X161Y130_BQ;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D3 = CLBLM_R_X89Y122_SLICE_X141Y122_BQ;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D4 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D5 = CLBLM_R_X89Y125_SLICE_X140Y125_DQ;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_D6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B5 = CLBLL_L_X102Y130_SLICE_X160Y130_CO6;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y122_SLICE_X141Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C1 = CLBLL_L_X102Y127_SLICE_X160Y127_BQ;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C2 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C3 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C4 = CLBLL_L_X102Y130_SLICE_X160Y130_B5Q;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_C5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A4 = CLBLM_R_X89Y122_SLICE_X140Y122_BO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A5 = CLBLM_R_X89Y126_SLICE_X141Y126_DO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A6 = CLBLM_L_X90Y121_SLICE_X142Y121_AQ;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B1 = CLBLM_R_X89Y122_SLICE_X140Y122_AQ;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B2 = CLBLM_R_X89Y122_SLICE_X140Y122_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B4 = CLBLM_R_X89Y122_SLICE_X140Y122_CQ;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B5 = CLBLM_R_X89Y122_SLICE_X140Y122_C5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_B6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D4 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D5 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X160Y129_D6 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C2 = CLBLM_R_X89Y122_SLICE_X140Y122_CQ;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C3 = CLBLM_R_X89Y122_SLICE_X140Y122_AQ;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C4 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C5 = 1'b1;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_C6 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A1 = CLBLM_R_X93Y129_SLICE_X146Y129_A5Q;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A3 = CLBLM_L_X92Y129_SLICE_X145Y129_BO6;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_A6 = CLBLM_R_X95Y131_SLICE_X150Y131_DO6;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_AX = CLBLM_L_X92Y129_SLICE_X145Y129_BO5;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_B1 = CLBLM_L_X92Y129_SLICE_X145Y129_AQ;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D1 = CLBLM_R_X89Y122_SLICE_X140Y122_C5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D2 = CLBLM_R_X89Y122_SLICE_X140Y122_AQ;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D3 = CLBLM_L_X92Y121_SLICE_X145Y121_C5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D4 = CLBLM_R_X89Y122_SLICE_X140Y122_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_D6 = CLBLM_R_X89Y122_SLICE_X140Y122_CQ;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A4 = CLBLL_L_X102Y130_SLICE_X161Y130_BQ;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A5 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A6 = CLBLM_R_X101Y128_SLICE_X158Y128_A5Q;
  assign CLBLM_R_X89Y122_SLICE_X140Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C2 = CLBLM_L_X92Y129_SLICE_X145Y129_CQ;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C3 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C4 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_C5 = CLBLM_L_X92Y129_SLICE_X145Y129_AQ;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_B6 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D1 = CLBLM_L_X92Y129_SLICE_X145Y129_C5Q;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D2 = CLBLM_L_X92Y129_SLICE_X145Y129_CQ;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D3 = CLBLM_L_X90Y128_SLICE_X143Y128_DQ;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D4 = CLBLM_L_X92Y129_SLICE_X145Y129_A5Q;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D5 = CLBLM_L_X92Y129_SLICE_X145Y129_AQ;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C1 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C5 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X145Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_C2 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A1 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A2 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A3 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A4 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A5 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_A6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D1 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D2 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D3 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D4 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D5 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B1 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B2 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B3 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B4 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B5 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_B6 = 1'b1;
  assign CLBLL_L_X102Y129_SLICE_X161Y129_D6 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C1 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C2 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C3 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C4 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C5 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_C6 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D1 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D2 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D3 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D4 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D5 = 1'b1;
  assign CLBLM_L_X92Y129_SLICE_X144Y129_D6 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A2 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A3 = CLBLM_R_X103Y121_SLICE_X163Y121_AQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A4 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A5 = CLBLM_R_X103Y120_SLICE_X163Y120_AQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_OLOGIC_X0Y81_T1 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B2 = CLBLM_R_X103Y122_SLICE_X163Y122_BQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B3 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B4 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B5 = CLBLM_R_X103Y121_SLICE_X163Y121_C5Q;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_B6 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C1 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C2 = CLBLM_R_X103Y121_SLICE_X163Y121_CQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C4 = CLBLM_R_X103Y122_SLICE_X163Y122_CQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C5 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_C6 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D1 = CLBLM_R_X103Y121_SLICE_X163Y121_C5Q;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D2 = CLBLM_R_X103Y121_SLICE_X163Y121_CQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D3 = CLBLM_R_X103Y122_SLICE_X163Y122_CQ;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D4 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D5 = CLBLM_R_X103Y121_SLICE_X163Y121_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y121_SLICE_X163Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A2 = CLBLM_R_X103Y121_SLICE_X162Y121_DO6;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A4 = CLBLM_R_X103Y120_SLICE_X162Y120_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_A6 = CLBLL_L_X100Y121_SLICE_X157Y121_DO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = 1'b0;
  assign LIOB33_X0Y123_IOB_X0Y124_O = 1'b0;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B2 = CLBLM_R_X103Y121_SLICE_X162Y121_BQ;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B3 = CLBLM_R_X103Y121_SLICE_X162Y121_AQ;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B4 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B5 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_B6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y123_T = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y124_T = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C1 = CLBLM_R_X103Y121_SLICE_X162Y121_BQ;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C2 = CLBLM_R_X103Y121_SLICE_X162Y121_AQ;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C3 = CLBLL_L_X102Y121_SLICE_X161Y121_A5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C5 = CLBLM_R_X103Y121_SLICE_X162Y121_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_C6 = CLBLM_R_X103Y120_SLICE_X162Y120_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D1 = CLBLM_R_X103Y121_SLICE_X162Y121_BQ;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D2 = CLBLM_R_X103Y121_SLICE_X162Y121_AQ;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D3 = CLBLL_L_X102Y121_SLICE_X161Y121_A5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D5 = CLBLM_R_X103Y121_SLICE_X162Y121_B5Q;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_D6 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A1 = CLBLM_R_X89Y123_SLICE_X141Y123_AQ;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A2 = CLBLM_L_X90Y121_SLICE_X143Y121_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A4 = CLBLM_L_X90Y123_SLICE_X142Y123_BQ;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A5 = CLBLM_R_X89Y122_SLICE_X140Y122_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_A6 = 1'b1;
  assign CLBLM_R_X103Y121_SLICE_X162Y121_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B1 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B2 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A2 = CLBLL_L_X102Y130_SLICE_X160Y130_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_B6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A4 = CLBLL_L_X102Y129_SLICE_X160Y129_AQ;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C1 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C2 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_A6 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_C6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B2 = CLBLL_L_X102Y130_SLICE_X160Y130_BQ;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B4 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B5 = CLBLL_L_X102Y129_SLICE_X160Y129_BQ;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_B6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C1 = CLBLL_L_X102Y129_SLICE_X160Y129_BQ;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C3 = CLBLL_L_X102Y129_SLICE_X160Y129_C5Q;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C4 = CLBLL_L_X102Y130_SLICE_X160Y130_BQ;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C5 = CLBLL_L_X102Y130_SLICE_X160Y130_B5Q;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_C6 = CLBLL_L_X102Y130_SLICE_X161Y130_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y123_SLICE_X141Y123_D3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D1 = CLBLL_L_X102Y129_SLICE_X160Y129_BQ;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D2 = CLBLL_L_X102Y129_SLICE_X160Y129_C5Q;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D3 = CLBLL_L_X102Y130_SLICE_X160Y130_BQ;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D5 = CLBLL_L_X102Y130_SLICE_X160Y130_B5Q;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_D6 = CLBLL_L_X100Y130_SLICE_X156Y130_AQ;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A1 = CLBLM_R_X89Y128_SLICE_X140Y128_DO6;
  assign CLBLL_L_X102Y130_SLICE_X160Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A4 = CLBLM_R_X89Y123_SLICE_X140Y123_BO6;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_A6 = CLBLM_R_X89Y124_SLICE_X140Y124_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_AX = CLBLM_R_X89Y123_SLICE_X140Y123_BO5;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B1 = CLBLM_R_X89Y123_SLICE_X140Y123_AQ;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B2 = CLBLM_R_X89Y123_SLICE_X140Y123_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B4 = CLBLM_R_X89Y123_SLICE_X140Y123_CQ;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B5 = CLBLM_R_X89Y123_SLICE_X140Y123_C5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_B6 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C2 = CLBLM_R_X89Y123_SLICE_X140Y123_CQ;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C3 = CLBLM_R_X89Y123_SLICE_X140Y123_AQ;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C4 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_C6 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A2 = CLBLL_L_X102Y130_SLICE_X161Y130_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D1 = CLBLM_R_X89Y123_SLICE_X140Y123_C5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D2 = CLBLM_R_X89Y123_SLICE_X140Y123_AQ;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D3 = CLBLM_L_X92Y123_SLICE_X144Y123_D5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D4 = CLBLM_R_X89Y123_SLICE_X140Y123_A5Q;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_D6 = CLBLM_R_X89Y123_SLICE_X140Y123_CQ;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A4 = CLBLL_L_X102Y134_SLICE_X160Y134_AQ;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_A5 = 1'b1;
  assign CLBLM_R_X89Y123_SLICE_X140Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B3 = CLBLL_L_X102Y129_SLICE_X160Y129_C5Q;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B4 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B5 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_B2 = CLBLM_R_X101Y135_SLICE_X159Y135_D5Q;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C1 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C4 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C5 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_C2 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D1 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D2 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D3 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D4 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D5 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_D6 = 1'b1;
  assign CLBLL_L_X102Y130_SLICE_X161Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A3 = CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A5 = CLBLM_R_X103Y122_SLICE_X162Y122_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B2 = CLBLM_R_X103Y122_SLICE_X163Y122_A5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B4 = CLBLL_L_X102Y121_SLICE_X160Y121_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B5 = CLBLM_R_X103Y122_SLICE_X163Y122_C5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C1 = CLBLL_L_X102Y122_SLICE_X161Y122_C5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C2 = CLBLM_R_X103Y122_SLICE_X162Y122_A5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C5 = CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = 1'b0;
  assign LIOB33_X0Y125_IOB_X0Y126_O = 1'b0;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y125_IOB_X0Y126_T = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_T = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D1 = CLBLM_R_X103Y122_SLICE_X162Y122_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D2 = CLBLM_R_X103Y123_SLICE_X163Y123_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D4 = CLBLM_R_X103Y122_SLICE_X163Y122_A5Q;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D6 = CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A2 = CLBLM_R_X103Y122_SLICE_X162Y122_B5Q;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A5 = CLBLM_R_X103Y123_SLICE_X163Y123_AQ;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B2 = CLBLM_R_X103Y122_SLICE_X162Y122_BQ;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B4 = CLBLM_R_X103Y123_SLICE_X162Y123_BQ;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C2 = CLBLL_L_X100Y122_SLICE_X157Y122_C5Q;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C3 = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C5 = CLBLM_R_X103Y121_SLICE_X163Y121_DO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C6 = CLBLL_L_X102Y121_SLICE_X161Y121_CQ;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D3 = CLBLM_R_X103Y122_SLICE_X162Y122_BQ;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D4 = CLBLM_R_X103Y122_SLICE_X162Y122_A5Q;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D5 = CLBLM_R_X103Y122_SLICE_X162Y122_B5Q;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D6 = CLBLM_R_X103Y123_SLICE_X162Y123_BQ;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A1 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A2 = CLBLM_R_X89Y124_SLICE_X141Y124_A5Q;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A4 = CLBLM_R_X89Y130_SLICE_X141Y130_AQ;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A5 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B2 = CLBLM_R_X89Y124_SLICE_X140Y124_BO6;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B5 = CLBLM_R_X89Y124_SLICE_X141Y124_A5Q;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A4 = CLBLM_R_X101Y131_SLICE_X159Y131_CQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_A6 = CLBLL_L_X102Y131_SLICE_X160Y131_CO6;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_B1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C2 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C3 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C4 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C5 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_C6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B2 = CLBLL_L_X102Y131_SLICE_X160Y131_BQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B3 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B4 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B5 = CLBLM_R_X101Y131_SLICE_X159Y131_BQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_B6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C1 = CLBLM_R_X101Y131_SLICE_X159Y131_BQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C2 = CLBLL_L_X102Y130_SLICE_X160Y130_A5Q;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C3 = CLBLL_L_X102Y131_SLICE_X160Y131_AQ;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D2 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D3 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D4 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D5 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_D6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C5 = CLBLL_L_X102Y131_SLICE_X160Y131_B5Q;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y124_SLICE_X141Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D1 = CLBLM_R_X101Y131_SLICE_X159Y131_BQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D2 = CLBLL_L_X102Y131_SLICE_X160Y131_AQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D3 = CLBLM_L_X98Y130_SLICE_X155Y130_DQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D4 = CLBLL_L_X102Y131_SLICE_X160Y131_BQ;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D5 = CLBLL_L_X102Y131_SLICE_X160Y131_B5Q;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y131_SLICE_X160Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A1 = CLBLM_L_X90Y125_SLICE_X143Y125_AQ;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A2 = CLBLM_R_X89Y124_SLICE_X140Y124_A5Q;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A4 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A5 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_A6 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B1 = CLBLM_R_X89Y125_SLICE_X140Y125_DQ;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B2 = CLBLM_R_X89Y124_SLICE_X140Y124_BQ;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B4 = CLBLM_R_X89Y124_SLICE_X141Y124_BQ;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B5 = CLBLM_R_X89Y122_SLICE_X141Y122_D5Q;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_B6 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A1 = CLBLM_L_X92Y131_SLICE_X145Y131_BO6;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C2 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C3 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C4 = CLBLM_R_X89Y121_SLICE_X140Y121_A5Q;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C5 = CLBLM_R_X89Y126_SLICE_X140Y126_B5Q;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_C6 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A3 = CLBLM_R_X93Y130_SLICE_X146Y130_BQ;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A5 = CLBLM_R_X97Y131_SLICE_X152Y131_CO6;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B5 = CLBLM_L_X92Y131_SLICE_X144Y131_AQ;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_B6 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D1 = CLBLM_R_X89Y122_SLICE_X141Y122_D5Q;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D2 = CLBLM_R_X89Y124_SLICE_X140Y124_CQ;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D3 = CLBLM_R_X89Y124_SLICE_X140Y124_BQ;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C1 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D4 = CLBLM_R_X89Y125_SLICE_X140Y125_DQ;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C2 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C3 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C4 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C5 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_C6 = 1'b1;
  assign CLBLM_R_X89Y124_SLICE_X140Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_B5 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D1 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D2 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D3 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D4 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D5 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_D6 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C4 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_C5 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X145Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D1 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D2 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A1 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A2 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D3 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D5 = 1'b1;
  assign CLBLL_L_X102Y131_SLICE_X161Y131_D6 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A3 = CLBLM_L_X92Y131_SLICE_X144Y131_AQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A5 = CLBLM_L_X92Y131_SLICE_X145Y131_AQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_A6 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B1 = CLBLM_L_X90Y131_SLICE_X142Y131_A5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B3 = CLBLM_L_X90Y128_SLICE_X143Y128_D5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B4 = CLBLM_L_X90Y130_SLICE_X142Y130_B5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B5 = CLBLM_L_X92Y131_SLICE_X144Y131_BQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_B6 = 1'b1;
  assign LIOI3_X0Y205_OLOGIC_X0Y206_D1 = 1'b0;
  assign LIOI3_X0Y205_OLOGIC_X0Y206_T1 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C2 = CLBLM_L_X92Y131_SLICE_X144Y131_CQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C3 = CLBLM_R_X89Y130_SLICE_X140Y130_AQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C4 = CLBLM_R_X89Y128_SLICE_X140Y128_A5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C5 = CLBLM_L_X92Y131_SLICE_X144Y131_B5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_C6 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y205_OLOGIC_X0Y205_D1 = 1'b0;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D1 = CLBLM_L_X92Y131_SLICE_X145Y131_AQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D2 = CLBLM_L_X92Y131_SLICE_X145Y131_A5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D3 = CLBLM_L_X92Y131_SLICE_X144Y131_AQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D4 = CLBLM_L_X92Y131_SLICE_X144Y131_A5Q;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D5 = CLBLM_L_X92Y131_SLICE_X144Y131_BQ;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_D1 = 1'b0;
  assign LIOI3_X0Y205_OLOGIC_X0Y205_T1 = 1'b1;
  assign CLBLM_L_X92Y131_SLICE_X144Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y83_OLOGIC_X0Y84_T1 = 1'b1;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_D1 = 1'b0;
  assign LIOB33_X0Y75_IOB_X0Y76_O = 1'b0;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_D1 = 1'b0;
  assign LIOI3_X0Y83_OLOGIC_X0Y83_T1 = 1'b1;
  assign LIOB33_X0Y75_IOB_X0Y75_O = 1'b0;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A1 = CLBLM_L_X92Y127_SLICE_X145Y127_BQ;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y208_T1 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOB33_X0Y127_IOB_X0Y128_O = 1'b0;
  assign LIOB33_X0Y127_IOB_X0Y127_O = 1'b0;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_A3 = CLBLM_L_X92Y127_SLICE_X145Y127_AQ;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_D1 = 1'b0;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = 1'b0;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A2 = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A3 = CLBLM_R_X103Y126_SLICE_X163Y126_DO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A5 = CLBLM_R_X103Y123_SLICE_X162Y123_AQ;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y127_IOB_X0Y127_T = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_T = 1'b1;
  assign LIOI3_TBYTESRC_X0Y207_OLOGIC_X0Y207_T1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B4 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B5 = CLBLM_R_X103Y122_SLICE_X163Y122_C5Q;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C1 = CLBLL_L_X102Y122_SLICE_X161Y122_C5Q;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C4 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C5 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y75_IOB_X0Y76_T = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D4 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B3 = CLBLM_R_X101Y112_SLICE_X159Y112_A5Q;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y75_IOB_X0Y75_T = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A2 = CLBLM_R_X103Y123_SLICE_X162Y123_A5Q;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A3 = CLBLM_R_X101Y123_SLICE_X159Y123_AQ;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A4 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A5 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B2 = CLBLM_R_X103Y123_SLICE_X163Y123_BO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B5 = CLBLM_R_X103Y123_SLICE_X162Y123_A5Q;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B6 = CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C1 = CLBLM_R_X101Y123_SLICE_X159Y123_AQ;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C2 = CLBLM_R_X103Y123_SLICE_X163Y123_CO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C3 = CLBLL_L_X102Y122_SLICE_X161Y122_DO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C5 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C3 = CLBLL_L_X102Y114_SLICE_X160Y114_BQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D5 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C4 = CLBLL_L_X102Y115_SLICE_X160Y115_B5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C4 = CLBLM_L_X92Y127_SLICE_X145Y127_AQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A2 = CLBLM_L_X92Y126_SLICE_X145Y126_DO6;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C5 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A4 = CLBLM_R_X89Y125_SLICE_X141Y125_BO6;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C5 = CLBLM_L_X92Y127_SLICE_X145Y127_B5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A5 = CLBLM_R_X89Y125_SLICE_X140Y125_AQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_AX = CLBLM_R_X89Y125_SLICE_X141Y125_BO5;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B1 = CLBLM_R_X89Y125_SLICE_X141Y125_AQ;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B2 = CLBLM_R_X89Y125_SLICE_X141Y125_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B4 = CLBLM_R_X89Y125_SLICE_X141Y125_CQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B5 = CLBLM_R_X89Y126_SLICE_X141Y126_C5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = 1'b0;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C2 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C3 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C4 = CLBLM_L_X90Y125_SLICE_X142Y125_AQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C5 = CLBLM_R_X89Y125_SLICE_X141Y125_AQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_C6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D1 = CLBLM_R_X89Y126_SLICE_X141Y126_C5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D2 = CLBLM_R_X89Y125_SLICE_X141Y125_CQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D3 = CLBLM_R_X89Y125_SLICE_X141Y125_AQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D4 = CLBLM_R_X89Y125_SLICE_X141Y125_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D5 = CLBLM_R_X89Y123_SLICE_X141Y123_AQ;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y125_SLICE_X141Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A1 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A2 = CLBLM_R_X89Y125_SLICE_X140Y125_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A4 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A5 = CLBLM_L_X90Y118_SLICE_X143Y118_AQ;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_A6 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B1 = CLBLM_R_X93Y126_SLICE_X147Y126_DO6;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D1 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B5 = CLBLM_R_X89Y125_SLICE_X140Y125_A5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_B6 = CLBLM_R_X89Y125_SLICE_X140Y125_CO6;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_BX = CLBLM_R_X89Y125_SLICE_X140Y125_CO5;
  assign CLBLM_L_X92Y127_SLICE_X145Y127_D2 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C2 = CLBLM_L_X90Y125_SLICE_X142Y125_AQ;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C3 = CLBLM_R_X89Y125_SLICE_X140Y125_BQ;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C4 = CLBLM_R_X89Y125_SLICE_X141Y125_C5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C5 = CLBLM_R_X89Y125_SLICE_X140Y125_B5Q;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_C6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_AX = CLBLM_L_X92Y132_SLICE_X145Y132_BO5;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_A1 = CLBLM_R_X95Y132_SLICE_X150Y132_DO6;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B1 = CLBLM_L_X92Y132_SLICE_X145Y132_AQ;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B2 = CLBLM_L_X92Y132_SLICE_X145Y132_A5Q;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B4 = CLBLM_L_X92Y132_SLICE_X145Y132_CQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B5 = CLBLM_L_X92Y132_SLICE_X145Y132_C5Q;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_B6 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D2 = CLBLM_R_X89Y128_SLICE_X140Y128_CQ;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D3 = CLBLM_R_X89Y124_SLICE_X141Y124_BQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C1 = CLBLM_L_X92Y132_SLICE_X145Y132_CQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C4 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C5 = CLBLM_L_X92Y132_SLICE_X145Y132_AQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_C6 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D4 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D5 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_D6 = 1'b1;
  assign CLBLM_R_X89Y125_SLICE_X140Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D1 = CLBLM_L_X92Y132_SLICE_X145Y132_C5Q;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D2 = CLBLM_L_X92Y132_SLICE_X145Y132_CQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D4 = CLBLM_L_X92Y132_SLICE_X145Y132_A5Q;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D5 = CLBLM_L_X92Y132_SLICE_X145Y132_AQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_D6 = CLBLM_L_X92Y131_SLICE_X144Y131_CQ;
  assign CLBLM_L_X92Y132_SLICE_X145Y132_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B2 = CLBLM_R_X101Y112_SLICE_X158Y112_B5Q;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A1 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A2 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A4 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A5 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_A6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B3 = CLBLL_L_X100Y111_SLICE_X156Y111_AQ;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B1 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B2 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B4 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B5 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_B6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_B6 = CLBLM_R_X101Y112_SLICE_X158Y112_CO6;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C1 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C2 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C4 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C5 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_C6 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_A4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = 1'b0;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D1 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D2 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D3 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D4 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D5 = 1'b1;
  assign CLBLM_L_X92Y132_SLICE_X144Y132_D6 = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = 1'b0;
  assign LIOB33_X0Y129_IOB_X0Y129_O = 1'b0;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_C6 = CLBLM_L_X98Y112_SLICE_X154Y112_BQ;
  assign LIOB33_X0Y129_IOB_X0Y130_T = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_T = 1'b1;
  assign CLBLL_L_X100Y112_SLICE_X156Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B5 = 1'b1;
  assign CLBLM_L_X92Y127_SLICE_X144Y127_B6 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A2 = CLBLL_L_X102Y124_SLICE_X160Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A4 = CLBLM_R_X103Y124_SLICE_X163Y124_DO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A5 = CLBLM_L_X98Y122_SLICE_X154Y122_DO6;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B2 = CLBLM_R_X103Y124_SLICE_X163Y124_BQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B3 = CLBLM_R_X103Y124_SLICE_X163Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B4 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B5 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_B6 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C2 = CLBLL_L_X102Y124_SLICE_X160Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C3 = CLBLL_L_X102Y124_SLICE_X160Y124_C5Q;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C4 = CLBLM_R_X103Y124_SLICE_X163Y124_BQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C5 = CLBLM_R_X103Y124_SLICE_X163Y124_B5Q;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_C6 = CLBLM_R_X103Y124_SLICE_X163Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D1 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D2 = CLBLM_R_X103Y124_SLICE_X163Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D3 = CLBLL_L_X102Y124_SLICE_X160Y124_C5Q;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D4 = CLBLM_R_X103Y124_SLICE_X163Y124_BQ;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D5 = CLBLM_R_X103Y124_SLICE_X163Y124_B5Q;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y124_SLICE_X163Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A2 = CLBLM_L_X98Y123_SLICE_X155Y123_DO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A4 = CLBLM_R_X103Y124_SLICE_X162Y124_DO6;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A5 = CLBLM_R_X103Y120_SLICE_X162Y120_AQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_A6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B2 = CLBLM_R_X103Y124_SLICE_X162Y124_BQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B3 = CLBLM_R_X103Y124_SLICE_X162Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B4 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B3 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B5 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_B6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B4 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C1 = CLBLM_R_X103Y120_SLICE_X162Y120_AQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C2 = CLBLM_R_X103Y124_SLICE_X162Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C3 = CLBLM_R_X103Y124_SLICE_X162Y124_BQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C5 = CLBLM_R_X103Y124_SLICE_X162Y124_B5Q;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_C6 = CLBLL_L_X102Y124_SLICE_X161Y124_A5Q;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C1 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D1 = 1'b1;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D2 = CLBLM_R_X103Y124_SLICE_X162Y124_AQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D3 = CLBLL_L_X102Y124_SLICE_X161Y124_A5Q;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D4 = CLBLM_R_X103Y124_SLICE_X162Y124_BQ;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D5 = CLBLM_R_X103Y124_SLICE_X162Y124_B5Q;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A4 = CLBLM_R_X89Y126_SLICE_X141Y126_BO6;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A5 = CLBLM_R_X93Y126_SLICE_X146Y126_DO6;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_A6 = CLBLM_R_X89Y127_SLICE_X141Y127_A5Q;
  assign CLBLM_R_X103Y124_SLICE_X162Y124_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_AX = CLBLM_R_X89Y126_SLICE_X141Y126_BO5;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B1 = CLBLM_R_X89Y128_SLICE_X141Y128_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B2 = CLBLM_R_X89Y126_SLICE_X141Y126_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B3 = CLBLM_R_X89Y126_SLICE_X141Y126_AQ;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B4 = CLBLM_R_X89Y126_SLICE_X141Y126_CQ;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_B6 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C2 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C3 = CLBLM_R_X89Y125_SLICE_X141Y125_CQ;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C4 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C5 = CLBLM_R_X89Y126_SLICE_X141Y126_AQ;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_C6 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C5 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C6 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D1 = CLBLM_R_X89Y123_SLICE_X141Y123_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D2 = CLBLM_R_X89Y128_SLICE_X141Y128_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D4 = CLBLM_R_X89Y126_SLICE_X141Y126_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D5 = CLBLM_R_X89Y126_SLICE_X141Y126_AQ;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_D6 = CLBLM_R_X89Y126_SLICE_X141Y126_CQ;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C3 = CLBLM_R_X93Y125_SLICE_X146Y125_AQ;
  assign CLBLM_R_X89Y126_SLICE_X141Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A2 = CLBLM_L_X90Y126_SLICE_X142Y126_AO6;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A5 = CLBLM_L_X90Y125_SLICE_X143Y125_AQ;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_A6 = CLBLM_R_X89Y130_SLICE_X140Y130_BO6;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B1 = CLBLM_L_X90Y126_SLICE_X142Y126_AQ;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B2 = CLBLM_R_X89Y123_SLICE_X140Y123_A5Q;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B4 = CLBLM_L_X90Y126_SLICE_X142Y126_C5Q;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B5 = CLBLM_R_X89Y126_SLICE_X140Y126_BQ;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_B6 = 1'b1;
  assign CLBLM_R_X93Y125_SLICE_X146Y125_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C1 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C2 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C3 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C4 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C5 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_C6 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D1 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D2 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D3 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D4 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D5 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_D6 = 1'b1;
  assign CLBLM_R_X89Y126_SLICE_X140Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X90Y129_SLICE_X142Y129_C3 = CLBLM_L_X90Y130_SLICE_X142Y130_BQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = 1'b0;
  assign LIOB33_X0Y131_IOB_X0Y131_O = 1'b0;
  assign LIOB33_X0Y131_IOB_X0Y132_T = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y131_T = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A1 = CLBLM_R_X103Y125_SLICE_X163Y125_DO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A3 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A5 = CLBLM_R_X103Y125_SLICE_X162Y125_AQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_A6 = CLBLM_R_X103Y126_SLICE_X163Y126_BO6;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B2 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B3 = CLBLM_R_X103Y125_SLICE_X163Y125_AQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B4 = CLBLM_R_X103Y125_SLICE_X162Y125_C5Q;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_B6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C2 = CLBLM_R_X103Y125_SLICE_X163Y125_CQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C4 = CLBLM_R_X103Y125_SLICE_X163Y125_BQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_C6 = 1'b1;
  assign LIOI3_X0Y209_OLOGIC_X0Y210_D1 = 1'b0;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y209_OLOGIC_X0Y210_T1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D1 = CLBLM_R_X103Y125_SLICE_X163Y125_C5Q;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D2 = CLBLM_R_X103Y125_SLICE_X163Y125_CQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D3 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D4 = CLBLM_R_X103Y125_SLICE_X163Y125_BQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D5 = CLBLM_R_X103Y125_SLICE_X163Y125_AQ;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y125_SLICE_X163Y125_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y209_OLOGIC_X0Y209_D1 = 1'b0;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A2 = CLBLM_R_X103Y125_SLICE_X162Y125_A5Q;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A3 = CLBLM_R_X103Y123_SLICE_X162Y123_AQ;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A4 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_A6 = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_D1 = 1'b0;
  assign LIOI3_X0Y209_OLOGIC_X0Y209_T1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B1 = CLBLM_R_X103Y126_SLICE_X163Y126_CO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B2 = CLBLM_R_X103Y125_SLICE_X162Y125_A5Q;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B3 = CLBLM_R_X103Y125_SLICE_X162Y125_DO6;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_B6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_T1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C1 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C2 = CLBLM_R_X103Y125_SLICE_X162Y125_CQ;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C4 = CLBLM_R_X103Y125_SLICE_X162Y125_BQ;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C5 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_C6 = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y85_D1 = 1'b0;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTESRC_X0Y219_OLOGIC_X0Y220_D1 = 1'b0;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D1 = CLBLM_R_X103Y125_SLICE_X162Y125_C5Q;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D2 = CLBLM_R_X103Y125_SLICE_X162Y125_CQ;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D3 = CLBLM_R_X103Y125_SLICE_X163Y125_B5Q;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A1 = CLBLM_R_X101Y136_SLICE_X158Y136_AQ;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A2 = CLBLL_L_X102Y134_SLICE_X160Y134_A5Q;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_A6 = 1'b1;
  assign CLBLM_R_X103Y125_SLICE_X162Y125_D4 = CLBLM_R_X103Y125_SLICE_X162Y125_BQ;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A2 = CLBLM_R_X89Y127_SLICE_X141Y127_A5Q;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A5 = CLBLM_R_X89Y125_SLICE_X140Y125_AQ;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_A6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B2 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B1 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B5 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B3 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_B4 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_B6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C1 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C2 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C3 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C5 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_C6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_C6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D1 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D2 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D4 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_D6 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y134_SLICE_X160Y134_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D6 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D3 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X141Y127_D5 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A3 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A5 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_A6 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B3 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B5 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_B6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A1 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A2 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C3 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C5 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_C6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_A6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B4 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_B6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C1 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D1 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D2 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D6 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_C6 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D4 = 1'b1;
  assign CLBLM_R_X89Y127_SLICE_X140Y127_D5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D1 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D2 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D3 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D4 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D5 = 1'b1;
  assign CLBLL_L_X102Y134_SLICE_X161Y134_D6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign LIOB33_X0Y133_IOB_X0Y133_O = 1'b0;
  assign LIOB33_X0Y133_IOB_X0Y134_T = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_T = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = 1'b0;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A2 = CLBLM_R_X103Y125_SLICE_X163Y125_B5Q;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A3 = CLBLM_R_X103Y122_SLICE_X163Y122_B5Q;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A4 = CLBLM_R_X103Y126_SLICE_X163Y126_AQ;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A5 = CLBLM_R_X103Y125_SLICE_X163Y125_C5Q;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_A6 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B2 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_B6 = CLBLM_R_X103Y126_SLICE_X163Y126_A5Q;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C2 = CLBLM_R_X103Y126_SLICE_X163Y126_AQ;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C5 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_C6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = 1'b0;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D4 = CLBLM_R_X103Y122_SLICE_X163Y122_B5Q;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_D6 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X163Y126_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A2 = CLBLL_L_X102Y126_SLICE_X161Y126_DQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A5 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_A6 = CLBLM_R_X103Y126_SLICE_X162Y126_CO6;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B2 = CLBLM_R_X103Y126_SLICE_X162Y126_BQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B3 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B4 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B5 = CLBLL_L_X102Y126_SLICE_X161Y126_BQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_B6 = 1'b1;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C1 = CLBLL_L_X102Y126_SLICE_X161Y126_BQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C2 = CLBLM_R_X103Y126_SLICE_X162Y126_AQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C3 = CLBLM_R_X103Y126_SLICE_X162Y126_BQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C4 = CLBLL_L_X102Y126_SLICE_X161Y126_A5Q;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C5 = CLBLM_R_X103Y126_SLICE_X162Y126_B5Q;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_C6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A2 = CLBLM_R_X101Y135_SLICE_X159Y135_D5Q;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A3 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A4 = CLBLL_L_X102Y135_SLICE_X160Y135_BO6;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D1 = CLBLL_L_X102Y126_SLICE_X161Y126_BQ;
  assign CLBLM_R_X103Y126_SLICE_X162Y126_D2 = CLBLM_R_X103Y126_SLICE_X162Y126_AQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B1 = CLBLM_R_X101Y135_SLICE_X158Y135_A5Q;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A1 = CLBLM_L_X90Y128_SLICE_X143Y128_CQ;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A2 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A4 = CLBLM_R_X89Y126_SLICE_X141Y126_CQ;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A5 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_A6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B3 = CLBLL_L_X102Y135_SLICE_X160Y135_AQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B4 = CLBLM_R_X101Y135_SLICE_X159Y135_AQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B5 = CLBLL_L_X102Y134_SLICE_X160Y134_AQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_B6 = CLBLM_R_X101Y135_SLICE_X158Y135_AQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C1 = CLBLL_L_X102Y136_SLICE_X160Y136_AQ;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B3 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C2 = CLBLL_L_X100Y134_SLICE_X156Y134_B5Q;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B5 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_B6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C3 = CLBLL_L_X102Y136_SLICE_X160Y136_BQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C4 = CLBLM_R_X101Y135_SLICE_X159Y135_BQ;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_C5 = CLBLL_L_X102Y136_SLICE_X160Y136_B5Q;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C1 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C2 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C3 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C4 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D1 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D2 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D3 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D4 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D5 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_D6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X160Y135_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_C6 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D1 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D2 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D3 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D4 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D5 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_D6 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X141Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A1 = CLBLM_R_X93Y130_SLICE_X147Y130_DO6;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A4 = CLBLM_R_X89Y128_SLICE_X140Y128_BO6;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A5 = CLBLM_R_X89Y130_SLICE_X141Y130_AQ;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_A6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_AX = CLBLM_R_X89Y128_SLICE_X140Y128_BO5;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A1 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A2 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A3 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B4 = CLBLM_R_X89Y128_SLICE_X140Y128_CQ;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B5 = CLBLM_R_X89Y125_SLICE_X140Y125_D5Q;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_B6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A4 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A5 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_A6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B1 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C2 = CLBLM_R_X89Y128_SLICE_X140Y128_AQ;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C3 = CLBLM_R_X89Y131_SLICE_X140Y131_AQ;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C4 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C5 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_C6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B2 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C1 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C2 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B5 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_B6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C3 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_C4 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D1 = CLBLM_R_X89Y125_SLICE_X140Y125_D5Q;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D2 = CLBLM_R_X89Y126_SLICE_X140Y126_B5Q;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D3 = CLBLM_R_X89Y128_SLICE_X140Y128_AQ;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D4 = CLBLM_R_X89Y128_SLICE_X140Y128_A5Q;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_D6 = CLBLM_R_X89Y128_SLICE_X140Y128_CQ;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D1 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D2 = 1'b1;
  assign CLBLM_R_X89Y128_SLICE_X140Y128_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D3 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D6 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D4 = 1'b1;
  assign CLBLL_L_X102Y135_SLICE_X161Y135_D5 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y135_T = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_T = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y79_T1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A4 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_A6 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B4 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_B6 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C4 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_C6 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D4 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X163Y127_D6 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A1 = CLBLL_L_X102Y127_SLICE_X161Y127_B5Q;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A2 = CLBLL_L_X102Y127_SLICE_X161Y127_CO6;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_A6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B4 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_B6 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C1 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C4 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C5 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_C6 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A4 = CLBLM_R_X101Y135_SLICE_X159Y135_C5Q;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_A6 = CLBLL_L_X102Y136_SLICE_X160Y136_CO6;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B1 = CLBLM_R_X101Y135_SLICE_X159Y135_BQ;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B3 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B5 = CLBLL_L_X102Y136_SLICE_X160Y136_BQ;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_B6 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D2 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D3 = 1'b1;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_D4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C1 = CLBLL_L_X102Y136_SLICE_X160Y136_BQ;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C2 = CLBLL_L_X102Y136_SLICE_X160Y136_AQ;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C3 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C4 = CLBLM_R_X101Y135_SLICE_X159Y135_BQ;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C5 = CLBLL_L_X102Y136_SLICE_X160Y136_B5Q;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_C6 = CLBLM_R_X101Y136_SLICE_X158Y136_AQ;
  assign CLBLM_R_X103Y127_SLICE_X162Y127_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D2 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D3 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D5 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_D6 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X160Y136_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y211_OLOGIC_X0Y212_D1 = 1'b0;
  assign LIOI3_X0Y211_OLOGIC_X0Y212_T1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A2 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A3 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A5 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_A6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = 1'b0;
  assign LIOB33_X0Y137_IOB_X0Y138_O = 1'b0;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B2 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B3 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B5 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_B6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_T = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y138_T = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_D1 = 1'b0;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C2 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C3 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C5 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_C6 = 1'b1;
  assign LIOI3_X0Y211_OLOGIC_X0Y211_T1 = 1'b1;
  assign RIOB33_X105Y59_IOB_X1Y59_O = 1'b0;
  assign RIOB33_X105Y59_IOB_X1Y60_O = 1'b0;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_T1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D1 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D2 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D3 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D4 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D5 = 1'b1;
  assign CLBLL_L_X102Y136_SLICE_X161Y136_D6 = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_D1 = 1'b0;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y232_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_D1 = 1'b0;
  assign RIOB33_X105Y59_IOB_X1Y60_T = 1'b1;
  assign RIOB33_X105Y59_IOB_X1Y59_T = 1'b1;
  assign LIOI3_TBYTESRC_X0Y231_OLOGIC_X0Y231_T1 = 1'b1;
  assign CLBLM_L_X98Y134_SLICE_X154Y134_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C3 = CLBLM_R_X101Y116_SLICE_X158Y116_DO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C5 = CLBLL_L_X102Y115_SLICE_X160Y115_DO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A2 = CLBLM_R_X89Y130_SLICE_X141Y130_A5Q;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A3 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A4 = CLBLM_L_X90Y130_SLICE_X142Y130_AQ;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A5 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_A6 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B1 = CLBLM_L_X92Y132_SLICE_X145Y132_DO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B2 = CLBLM_R_X89Y130_SLICE_X141Y130_A5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C4 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B3 = CLBLM_R_X89Y130_SLICE_X140Y130_AO6;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_B6 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOB33_X0Y221_IOB_X0Y222_O = 1'b0;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C1 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C2 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_C6 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C4 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C5 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C3 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_C6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y139_O = 1'b0;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y139_IOB_X0Y140_O = 1'b0;
  assign LIOB33_X0Y221_IOB_X0Y221_O = 1'b0;
  assign LIOB33_X0Y139_IOB_X0Y140_T = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D1 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D2 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D3 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D4 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D5 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_D6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y139_T = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X141Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A1 = CLBLM_R_X89Y130_SLICE_X141Y130_BQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A2 = CLBLM_R_X89Y131_SLICE_X140Y131_AQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A3 = CLBLM_R_X89Y130_SLICE_X140Y130_AQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A5 = CLBLM_R_X89Y128_SLICE_X140Y128_C5Q;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_A6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D3 = CLBLL_L_X102Y115_SLICE_X160Y115_BQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B1 = CLBLM_R_X89Y131_SLICE_X140Y131_AQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B3 = CLBLM_R_X89Y130_SLICE_X140Y130_AQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B4 = CLBLM_R_X89Y130_SLICE_X141Y130_BQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B5 = CLBLM_R_X89Y128_SLICE_X140Y128_C5Q;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_B6 = CLBLM_R_X89Y126_SLICE_X140Y126_BQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C1 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C2 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C3 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C4 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C5 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_C6 = 1'b1;
  assign LIOB33_X0Y221_IOB_X0Y222_T = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D3 = CLBLM_L_X92Y128_SLICE_X145Y128_CQ;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D1 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D2 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D3 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D4 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D5 = 1'b1;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_D6 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D4 = CLBLM_L_X92Y128_SLICE_X145Y128_A5Q;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D5 = CLBLM_L_X92Y128_SLICE_X145Y128_AQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X89Y130_SLICE_X140Y130_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X92Y128_SLICE_X145Y128_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B2 = CLBLL_L_X100Y113_SLICE_X156Y113_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b0;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B3 = CLBLL_L_X100Y113_SLICE_X156Y113_AQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C4 = CLBLL_L_X100Y112_SLICE_X157Y112_A5Q;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_A6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C5 = CLBLL_L_X100Y113_SLICE_X156Y113_B5Q;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X92Y128_SLICE_X144Y128_B1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b0;
  assign LIOI3_X0Y203_OLOGIC_X0Y204_T1 = 1'b1;
  assign CLBLM_L_X90Y130_SLICE_X143Y130_D5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign LIOI3_X0Y203_OLOGIC_X0Y203_D1 = 1'b0;
  assign LIOB33_X0Y141_IOB_X0Y142_O = 1'b0;
  assign LIOB33_X0Y141_IOB_X0Y141_O = 1'b0;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_A6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y141_T = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_T = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_B6 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_C6 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X141Y131_D6 = 1'b1;
  assign LIOI3_X0Y203_OLOGIC_X0Y203_T1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A1 = CLBLM_L_X90Y131_SLICE_X142Y131_CQ;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A5 = CLBLM_R_X89Y130_SLICE_X141Y130_BQ;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_A6 = 1'b1;
  assign CLBLM_L_X94Y122_SLICE_X149Y122_C2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B6 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_B5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_C6 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C6 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D1 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D2 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D3 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D4 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D5 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_D6 = 1'b1;
  assign CLBLM_R_X89Y131_SLICE_X140Y131_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y215_OLOGIC_X0Y216_D1 = 1'b0;
  assign LIOI3_X0Y215_OLOGIC_X0Y216_T1 = 1'b1;
  assign LIOI3_X0Y215_OLOGIC_X0Y215_D1 = 1'b0;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_D1 = 1'b0;
  assign LIOI3_X0Y215_OLOGIC_X0Y215_T1 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_T1 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_D1 = 1'b0;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y244_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y243_OLOGIC_X0Y243_T1 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = 1'b0;
  assign LIOB33_X0Y143_IOB_X0Y143_T = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOB33_SING_X105Y50_IOB_X1Y50_O = 1'b0;
  assign RIOB33_SING_X105Y50_IOB_X1Y50_T = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = 1'b0;
  assign LIOB33_X0Y145_IOB_X0Y145_O = 1'b0;
  assign RIOB33_SING_X105Y99_IOB_X1Y99_O = CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  assign LIOB33_X0Y145_IOB_X0Y146_T = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y145_T = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A2 = CLBLM_R_X97Y111_SLICE_X153Y111_A5Q;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A3 = CLBLM_R_X97Y112_SLICE_X153Y112_AQ;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A4 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A5 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_A6 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B1 = CLBLM_L_X98Y111_SLICE_X154Y111_CO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B2 = CLBLL_L_X100Y111_SLICE_X157Y111_B5Q;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B3 = CLBLM_R_X97Y112_SLICE_X153Y112_AQ;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B4 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B5 = CLBLM_L_X94Y111_SLICE_X149Y111_DO6;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_B6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C1 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C2 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C3 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C4 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C5 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_C6 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D1 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D2 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D3 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D4 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D5 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_D6 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X153Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A2 = CLBLM_R_X97Y112_SLICE_X152Y112_A5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A3 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A4 = CLBLM_R_X95Y111_SLICE_X150Y111_B5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A5 = CLBLM_R_X97Y111_SLICE_X152Y111_CO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_A6 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B2 = CLBLM_R_X97Y111_SLICE_X152Y111_BQ;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B3 = CLBLM_R_X97Y111_SLICE_X152Y111_AQ;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B4 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B5 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_B6 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C2 = CLBLM_R_X97Y111_SLICE_X153Y111_A5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C3 = CLBLM_R_X95Y111_SLICE_X150Y111_DO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C5 = CLBLM_R_X97Y111_SLICE_X152Y111_DO6;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_C6 = CLBLM_L_X98Y111_SLICE_X155Y111_A5Q;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_D1 = 1'b0;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D1 = CLBLM_R_X97Y111_SLICE_X152Y111_BQ;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D2 = CLBLM_R_X97Y111_SLICE_X152Y111_AQ;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D3 = CLBLM_L_X98Y111_SLICE_X155Y111_B5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D4 = 1'b1;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D5 = CLBLM_R_X97Y111_SLICE_X152Y111_B5Q;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_D6 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X97Y111_SLICE_X152Y111_SR = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_O = 1'b0;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_T1 = 1'b1;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_T = 1'b1;
endmodule
