module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD
  );
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_F7AMUX_O;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CLK;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_SR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_F7BMUX_O;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_SR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_SR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_SR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_SR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5d00ff000000cc)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc400ccf8c400cc)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0004040000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500aafaaaff)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X2Y110_SLICE_X1Y110_MUXF7A (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_BO6),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.O(CLBLL_L_X2Y110_SLICE_X1Y110_F7AMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacafafa0a0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h303000003c0c3232)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50d05054107034a4)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cc00000033cc)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a880080fffbf5ff)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88fcfcbb883030)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400a680110055cc)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X2Y111_SLICE_X1Y111_MUXF7A (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O(CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c200000002)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000a00000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222244444444)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03000000ff000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y101_IOB_X0Y101_I),
.D(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.Q(CLBLL_L_X2Y112_SLICE_X1Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ecc4ece0a404e04)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a8aa8820202200)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_F7AMUX_O),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_F7AMUX_O),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h030e000e03020002)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e080800000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X2Y112_SLICE_X1Y112_MUXF7A (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_BO6),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.O(CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200331122002200)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0000c000220000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000030)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033000020002000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLL_L_X2Y113_SLICE_X0Y113_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffbefffdff7d)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffebffffffffff)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33aaaafc30)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2301230122002200)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y114_SLICE_X0Y114_BO6),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000002000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000400000a840)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aac0aa00000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdecfdec31203120)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.I3(CLBLL_L_X2Y114_SLICE_X1Y114_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y114_SLICE_X1Y114_BO6),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff0ccefcff0ccf)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3060101000005500)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a080808080)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000303400000004)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X2Y115_SLICE_X0Y115_MUXF7A (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.O(CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h037f030000000000)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0cceeeec0ccee)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff77ab55ab)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5cdf18df5fdf1bdf)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf0fffff4f0fffff)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y111_SLICE_X4Y111_MUXF7A (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.O(CLBLL_L_X4Y111_SLICE_X4Y111_F7AMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y111_SLICE_X4Y111_MUXF7B (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.O(CLBLL_L_X4Y111_SLICE_X4Y111_F7BMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y101_IOB_X0Y101_I),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y101_IOB_X0Y101_I),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h17c357c300b000b0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h43100310000c000c)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa3aca000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_F7AMUX_O),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_F7BMUX_O),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa88a0000088a0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_F7AMUX_O),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ffd0ffff000f000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fb30c803fb70c84)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222227250ffff)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa55aa7daa7d)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y112_SLICE_X5Y112_MUXF7A (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.O(CLBLL_L_X4Y112_SLICE_X5Y112_F7AMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hec0ce000cc0cc000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f0d43014e0c4200)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0a0a0505005f00)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y109_SLICE_X2Y109_MUXF7A (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.O(CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y101_IOB_X0Y101_I),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8fafa44004400)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb080b080b0b08080)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_F7AMUX_O),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000200000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2aaa0aaaaaaaaaaa)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y109_SLICE_X3Y109_MUXF7A (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.O(CLBLM_R_X3Y109_SLICE_X3Y109_F7AMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdfdf13ffffff33)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb3ececff7f2020)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffefffeffceffc)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h550055335500ff00)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y110_SLICE_X2Y110_MUXF7A (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.O(CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccafafa0a0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333dfff3333ffff)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000808000cc80cc)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc1c0c0c002030303)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y101_IOB_X0Y101_I),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0ffccf3c03300)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf080fffff0f00000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0343d2d200008c8c)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000acac0000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ffff3333)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54ae04ae04)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000008008000)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000054550000ab)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000000ff000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a000005f5fffff)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h23ff230033773377)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd5d555577777777)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y112_SLICE_X2Y112_MUXF7A (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.O(CLBLM_R_X3Y112_SLICE_X2Y112_F7AMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y101_IOB_X0Y101_I),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h333371f12020b0b0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000e020e020)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_F7AMUX_O),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h05bd05bd001d00bd)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f830f830f430f4)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y112_SLICE_X3Y112_MUXF7A (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.O(CLBLM_R_X3Y112_SLICE_X3Y112_F7AMUX_O),
.S(CLBLM_R_X3Y111_SLICE_X2Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5a0f5a0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefffbffffeeee)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1a0500001a050001)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80800b8b80800888)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fffff0f0f)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa3afa3aca0aca0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f303a3fffffff3)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001303030300101)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00040c0c00040000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0fafacfc00a0a)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330000aaaa0000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc0000c4cc)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000008833000088)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h333322e2000022e2)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aa0a0050f0a0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y114_SLICE_X3Y114_MUXF7A (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.O(CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4455440050555000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_AO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f8f0a0200000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_CQ),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X3Y115_SLICE_X2Y115_MUXF7A (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.O(CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O),
.S(CLBLM_R_X3Y109_SLICE_X3Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_DO6),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_DO6),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_DO6),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X1Y114_DO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_AMUX = CLBLL_L_X2Y110_SLICE_X1Y110_F7AMUX_O;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_AMUX = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_BMUX = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_AMUX = CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_CMUX = CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_DMUX = CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_AMUX = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_BMUX = CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_AMUX = CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_DMUX = CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_AMUX = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_CMUX = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_AMUX = CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_BMUX = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_F7AMUX_O;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CMUX = CLBLL_L_X4Y111_SLICE_X4Y111_F7BMUX_O;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_AMUX = CLBLL_L_X4Y112_SLICE_X5Y112_F7AMUX_O;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CMUX = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AMUX = CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CMUX = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_AMUX = CLBLM_R_X3Y109_SLICE_X3Y109_F7AMUX_O;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_CMUX = CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_BMUX = CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_DMUX = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_BMUX = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AMUX = CLBLM_R_X3Y112_SLICE_X2Y112_F7AMUX_O;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_CMUX = CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_DMUX = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_F7AMUX_O;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_BMUX = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AMUX = CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AMUX = CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_SR = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_AX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = CLBLM_R_X3Y112_SLICE_X2Y112_F7AMUX_O;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = CLBLL_L_X2Y110_SLICE_X1Y110_F7AMUX_O;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_SR = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_SR = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_F7AMUX_O;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_F7AMUX_O;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLM_R_X3Y109_SLICE_X2Y109_F7AMUX_O;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_F7AMUX_O;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X3Y114_SLICE_X3Y114_F7AMUX_O;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_SR = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLL_L_X2Y111_SLICE_X1Y111_F7AMUX_O;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_AX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = CLBLM_R_X3Y109_SLICE_X3Y109_F7AMUX_O;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X2Y112_SLICE_X1Y112_F7AMUX_O;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_SR = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AX = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X3Y115_SLICE_X2Y115_F7AMUX_O;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_F7BMUX_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_AX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLL_L_X2Y112_SLICE_X1Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AX = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_F7AMUX_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_F7AMUX_O;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
endmodule
