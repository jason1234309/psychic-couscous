module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  input LIOB33_X0Y129_IOB_X0Y129_IPAD,
  input LIOB33_X0Y129_IOB_X0Y130_IPAD,
  input LIOB33_X0Y131_IOB_X0Y131_IPAD,
  input LIOB33_X0Y131_IOB_X0Y132_IPAD,
  input LIOB33_X0Y133_IOB_X0Y133_IPAD,
  input LIOB33_X0Y133_IOB_X0Y134_IPAD,
  input LIOB33_X0Y135_IOB_X0Y135_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output RIOB33_SING_X105Y100_IOB_X1Y100_OPAD,
  output RIOB33_X105Y101_IOB_X1Y101_OPAD,
  output RIOB33_X105Y101_IOB_X1Y102_OPAD,
  output RIOB33_X105Y103_IOB_X1Y103_OPAD,
  output RIOB33_X105Y103_IOB_X1Y104_OPAD,
  output RIOB33_X105Y105_IOB_X1Y105_OPAD,
  output RIOB33_X105Y105_IOB_X1Y106_OPAD,
  output RIOB33_X105Y107_IOB_X1Y107_OPAD,
  output RIOB33_X105Y107_IOB_X1Y108_OPAD,
  output RIOB33_X105Y109_IOB_X1Y109_OPAD,
  output RIOB33_X105Y109_IOB_X1Y110_OPAD,
  output RIOB33_X105Y111_IOB_X1Y111_OPAD,
  output RIOB33_X105Y111_IOB_X1Y112_OPAD,
  output RIOB33_X105Y113_IOB_X1Y113_OPAD,
  output RIOB33_X105Y113_IOB_X1Y114_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD
  );
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CLK;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_SR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CLK;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5Q;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_SR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AQ;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BQ;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CLK;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_SR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CLK;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_SR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CLK;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_SR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CLK;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_SR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5Q;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CLK;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_SR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_SR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_SR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_SR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_SR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5Q;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_SR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_SR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_SR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_SR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_SR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_SR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_SR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_SR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5Q;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_SR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_SR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5Q;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_SR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_SR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5Q;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_SR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_AO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_AO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_A_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_BO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_BO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_B_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_CO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_CO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_C_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_DO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_DO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X78Y113_D_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_AO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_AO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_A_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_BO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_BO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_B_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_CO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_CO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_C_XOR;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D1;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D2;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D3;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D4;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_DO5;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_DO6;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D_CY;
  wire [0:0] CLBLL_L_X52Y113_SLICE_X79Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_SR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5Q;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5Q;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_SR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CLK;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_SR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5Q;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CLK;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_SR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_SR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_SR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5Q;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_SR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_SR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_SR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5Q;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_SR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5Q;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_SR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_SR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5Q;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5Q;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_SR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_SR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5Q;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CLK;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_SR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5Q;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CLK;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_SR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5Q;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CLK;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_SR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CLK;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_SR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_SR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_SR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_SR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_SR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_SR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_SR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_SR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_SR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_SR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_SR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_SR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_SR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_SR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_SR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_SR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_SR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_SR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_O;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_O;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_O;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_O;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_O;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_O;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_O;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1;
  wire [0:0] RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y101_TQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_D1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_OQ;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_T1;
  wire [0:0] RIOI3_X105Y101_OLOGIC_X1Y102_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y103_TQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_D1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_OQ;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_T1;
  wire [0:0] RIOI3_X105Y103_OLOGIC_X1Y104_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y105_TQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_D1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_OQ;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_T1;
  wire [0:0] RIOI3_X105Y105_OLOGIC_X1Y106_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y109_TQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_D1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_OQ;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_T1;
  wire [0:0] RIOI3_X105Y109_OLOGIC_X1Y110_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y111_TQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_D1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_OQ;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_T1;
  wire [0:0] RIOI3_X105Y111_OLOGIC_X1Y112_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X0Y115_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X0Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f0aafa33f0aafa)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f222f222f222f22)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0a0a0ffececec)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y129_IOB_X0Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_C5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_D5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8ff88f8f88888)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(LIOB33_X0Y129_IOB_X0Y129_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0a0a0ffececec)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(LIOB33_X0Y129_IOB_X0Y129_I),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaaaeaeaeae)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0a0a0a0a)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff55ff55)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y123_IOB_X0Y124_I),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h050f050f55ff55ff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(1'b1),
.I2(LIOB33_X0Y129_IOB_X0Y129_I),
.I3(LIOB33_X0Y131_IOB_X0Y131_I),
.I4(1'b1),
.I5(LIOB33_X0Y121_IOB_X0Y121_I),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96699669fff0ffff)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.I2(LIOB33_X0Y119_IOB_X0Y119_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_X0Y129_IOB_X0Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heccfcccfcccfcccf)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(LIOB33_X0Y129_IOB_X0Y129_I),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7ff070ff7f0000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_DO6),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeed5aa5eddea55a)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I2(LIOB33_X0Y119_IOB_X0Y119_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffffffafffa)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I2(LIOB33_X0Y119_IOB_X0Y119_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_A5Q),
.Q(CLBLL_L_X2Y120_SLICE_X1Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y120_SLICE_X1Y120_AQ),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y120_SLICE_X1Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff5fff5f)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y129_IOB_X0Y129_I),
.I3(LIOB33_X0Y119_IOB_X0Y120_I),
.I4(1'b1),
.I5(LIOB33_X0Y119_IOB_X0Y119_I),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffffff)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y119_IOB_X0Y119_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I5(LIOB33_X0Y119_IOB_X0Y120_I),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y119_IOB_X0Y120_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y119_IOB_X0Y119_I),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(LIOB33_X0Y121_IOB_X0Y121_I),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y121_SLICE_X0Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y121_SLICE_X0Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafffffffff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y121_IOB_X0Y122_I),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c00100010)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffdff000a000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(LIOB33_X0Y121_IOB_X0Y122_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55000c00fff3aaff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I3(LIOB33_X0Y123_IOB_X0Y123_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y121_SLICE_X1Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0fffffff4fff)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(LIOB33_X0Y121_IOB_X0Y121_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fe00eeffffffff)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(LIOB33_X0Y127_IOB_X0Y127_I),
.I1(LIOB33_X0Y127_IOB_X0Y128_I),
.I2(LIOB33_X0Y129_IOB_X0Y130_I),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0f0f0fcc00cc00)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_A5Q),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X0Y122_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_B5Q),
.I4(LIOB33_X0Y131_IOB_X0Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbf88888888)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(LIOB33_X0Y121_IOB_X0Y122_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y122_SLICE_X0Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y122_SLICE_X0Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_D5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0c0c0c0c)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_BQ),
.I2(LIOB33_X0Y133_IOB_X0Y134_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_CQ),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3230000055ff55ff)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_B5Q),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I2(LIOB33_X0Y135_IOB_X0Y135_I),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03fc30cf03fc30)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55665555)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdf)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcf0303cffc0330)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0f0f0f3c)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000101fefe)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y103_IOB_X0Y104_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafac8c8c8c8)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5703ffff5703ffff)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_B5Q),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff44ff50ff50)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5500ffff4444)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y101_IOB_X0Y101_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccff66999966)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00200000fffbffff)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f7b3f7b55ff0000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f0f5f0f5f0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00ff00f0ff0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_CQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_DQ),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55a5aa55aa5a55a)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_C5Q),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_A5Q),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696696969699696)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_AQ),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_D5Q),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h08080088eeeeffff)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_CQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7f7fffff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_CQ),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I5(LIOB33_X0Y125_IOB_X0Y126_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010003000100)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200070)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbffcbfcfffcfff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_DQ),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a8fcfca8a8fcfc)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0357ffff0357ffff)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h220a000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I1(CLBLL_L_X2Y115_SLICE_X0Y115_CQ),
.I2(CLBLL_L_X2Y115_SLICE_X0Y115_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00040c0403000300)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_A5Q),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I4(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf8c8c8c8c)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X0Y115_AQ),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_A5Q),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055ffff3377ffff)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_CQ),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaa8aa)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00010031cfffcfff)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04000000c4000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdffffffdddf)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800f8f070f0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010011000100)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005300000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_DQ),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0ff0000000f)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000400000004000c)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_A5Q),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbffff7777ffff)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h12303030ffffefff)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff8fffa)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888888888cc8)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f00ff000c005d)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdfff0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000020)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff05370505)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_A5Q),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_A5Q),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcf6f6f3f6f)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3233223300000000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000000020000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3ffcfcfcfc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeffaaefeaffaa)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff0fcf0fd)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_A5Q),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000cc50dc)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8a8f0a07777ffff)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_D5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040004080800000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5757575700570000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550055000c0000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f2fafa)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000e0eff00)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff10ff00)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_A5Q),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000000)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffff00000010)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fff40000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0353005003030000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_A5Q),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000008000000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffffff)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005050cc00cc00)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8a8ffffa8ff)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_CO6),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_CQ),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X78Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X78Y113_DO5),
.O6(CLBLL_L_X52Y113_SLICE_X78Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X78Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X78Y113_CO5),
.O6(CLBLL_L_X52Y113_SLICE_X78Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X78Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X78Y113_BO5),
.O6(CLBLL_L_X52Y113_SLICE_X78Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X52Y113_SLICE_X78Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X78Y113_AO5),
.O6(CLBLL_L_X52Y113_SLICE_X78Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X79Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X79Y113_DO5),
.O6(CLBLL_L_X52Y113_SLICE_X79Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X79Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X79Y113_CO5),
.O6(CLBLL_L_X52Y113_SLICE_X79Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X79Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X79Y113_BO5),
.O6(CLBLL_L_X52Y113_SLICE_X79Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y113_SLICE_X79Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y113_SLICE_X79Y113_AO5),
.O6(CLBLL_L_X52Y113_SLICE_X79Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y105_IOB_X0Y106_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y107_IOB_X0Y108_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff7ffff)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0aff0a0a0aff0a)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff00ff55550000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ff44ff44444444)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I4(1'b1),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_C5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffecececffa0a0a0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefaaafcccf000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y129_IOB_X0Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf0cc00fefaeeaa)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e4eff44e4e4ff44)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22f2f222eef2f2)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y103_IOB_X0Y103_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y101_IOB_X0Y102_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff03330fff03330)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_A5Q),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0357ffff00ff00ff)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeccaa00fefcfaf0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y129_IOB_X0Y129_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I3(LIOB33_X0Y131_IOB_X0Y131_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y105_IOB_X0Y105_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y107_IOB_X0Y107_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5a9aaa9aa)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0e1f0e1)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ffcfcfc00)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I4(CLBLL_L_X2Y115_SLICE_X1Y115_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_BQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(LIOB33_X0Y109_IOB_X0Y109_I),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccaa88aa88)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeeee00ee00)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_DQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff0aff0affffff)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_C5Q),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f1fffff1111ffff)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_D5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ffbbbb00ccaaaa)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff96696996)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DQ),
.I3(CLBLL_L_X2Y115_SLICE_X0Y115_CQ),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heee0fff00f0f0f0f)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_A5Q),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_BQ),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0c0c0ffeaeaea)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffa000ffff0000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_B5Q),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaaacaaaaaaaaaaa)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_C5Q),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_CQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55557777ff55ff77)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_CQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_A5Q),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_C5Q),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_CQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330303cc001111)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I1(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DQ),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_A5Q),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9fbffffdfffdfff)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(LIOB33_X0Y121_IOB_X0Y121_I),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fccf0ccaaeeaaee)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfaf0eeccaa00)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y131_IOB_X0Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007700ff88ff00ff)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_D5Q),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I5(CLBLL_L_X2Y115_SLICE_X0Y115_BQ),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f7f0f3f5f7f0f3)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_DO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000200000002a)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_CQ),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001002300)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbf1fff5fffff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(LIOB33_X0Y121_IOB_X0Y121_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(LIOB33_X0Y123_IOB_X0Y124_I),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h35350000fafaffff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(1'b1),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h153f153f030f33ff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(LIOB33_X0Y123_IOB_X0Y123_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y123_IOB_X0Y124_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000a000008080)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y121_IOB_X0Y121_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h057f7fff5f7f7fff)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(LIOB33_X0Y123_IOB_X0Y124_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y123_IOB_X0Y123_I),
.I5(LIOB33_X0Y121_IOB_X0Y121_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h12003000efffffff)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaeaeaeaea)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I1(LIOB33_X0Y129_IOB_X0Y129_I),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_DO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc000ffffc000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_A5Q),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000010000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007700ff0000ffff)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_BQ),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f003f0000007fff)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_BQ),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33733777ccdccddd)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(LIOB33_X0Y123_IOB_X0Y123_I),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(LIOB33_X0Y123_IOB_X0Y124_I),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa88880a000800)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafa0f3f5a7b)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff00000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_B5Q),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLL_L_X2Y122_SLICE_X0Y122_AQ),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffaaffea)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I4(LIOB33_X0Y133_IOB_X0Y133_I),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h080000000f000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_B5Q),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_A5Q),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_AQ),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000030301010)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000030331011)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1333333333333333)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I1(LIOB33_X0Y135_IOB_X0Y135_I),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_A5Q),
.I5(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020004000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffffffffffff)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_BQ),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_A5Q),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf0f0faaaa0000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(1'b0),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_A5Q),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_BQ),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc800c000fa00f000)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_A5Q),
.I2(LIOB33_X0Y135_IOB_X0Y135_I),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_D5Q),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_B5Q),
.I5(CLBLL_L_X2Y122_SLICE_X0Y122_AQ),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff0f0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_A5Q),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y122_SLICE_X3Y122_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y122_SLICE_X3Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fe01ff00fe01)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_A5Q),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X3Y123_SLICE_X3Y123_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_DQ),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee00eee0e000e0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f6f6f999666699)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f69966f6f96699)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77777777ffffffff)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_B5Q),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fcc0caa0a8808)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_B5Q),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55aa55a5aa55aa5)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996699666699)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_A5Q),
.I5(CLBLL_L_X2Y115_SLICE_X1Y115_B5Q),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hebc3be3cbe3cebc3)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I2(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cccc33cc3333cc)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f00cccc0c00)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ccaaaa0088)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f1f1fffffefef)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0fff1fef)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300f3f0f3f0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0fff5f5f5fff)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeee0e000ee00e0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_DQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5affa5a5a5)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_A5Q),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f333f300f000f0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222f2f22222f2f2)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0acececece)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c0a080ffccaa88)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CQ),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f333f300f000f0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff44f040f040)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fcc0caa0a8808)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_DQ),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbfbfbfffffffff)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff333300ff0000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0f3f0a2a0a2a0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_B5Q),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000100ff00fe00)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c480044cc88)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeff00000400)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcf0fcf00cc00cc)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22222222ff22ff22)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00cfcccfcc)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fbfd0000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee2eeeeeffffff3f)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffff22202222)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ffffff6ffff6)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h006c00c0006000c0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_B5Q),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BQ),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999aa999999aaaa)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000200)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffedfffffffffff)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_A5Q),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1313000001320000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_A5Q),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccffffffff)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_D5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0000001e00)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h400000000000ffff)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DQ),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_D5Q),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffffff)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000444400044440)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_CQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf0f088ff88ff)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66666666f9f99999)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_A5Q),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1eff1eff11111111)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_B5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff77ffff3f0fcf)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_B5Q),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cccccc44444488)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ffb0ffffffffff)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A5_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3ececb3ecb3b3ec)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_A5Q),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_B5Q),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fc33c3cc3)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_A5Q),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_B5Q),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.PRE(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y129_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y129_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y130_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y130_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y131_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y131_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y132_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y132_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y133_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y134_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y135_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y101_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.O(RIOB33_X105Y101_IOB_X1Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y101_IOB_X1Y102_OBUF (
.I(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.O(RIOB33_X105Y101_IOB_X1Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y103_OBUF (
.I(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.O(RIOB33_X105Y103_IOB_X1Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y103_IOB_X1Y104_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.O(RIOB33_X105Y103_IOB_X1Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y105_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.O(RIOB33_X105Y105_IOB_X1Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y105_IOB_X1Y106_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.O(RIOB33_X105Y105_IOB_X1Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y107_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.O(RIOB33_X105Y107_IOB_X1Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y107_IOB_X1Y108_OBUF (
.I(1'b1),
.O(RIOB33_X105Y107_IOB_X1Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y109_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.O(RIOB33_X105Y109_IOB_X1Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y109_IOB_X1Y110_OBUF (
.I(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.O(RIOB33_X105Y109_IOB_X1Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y111_OBUF (
.I(1'b1),
.O(RIOB33_X105Y111_IOB_X1Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y111_IOB_X1Y112_OBUF (
.I(CLBLL_L_X52Y113_SLICE_X78Y113_AO6),
.O(RIOB33_X105Y111_IOB_X1Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y113_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O(RIOB33_X105Y113_IOB_X1Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y113_IOB_X1Y114_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.O(RIOB33_X105Y113_IOB_X1Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y100_IOB_X1Y100_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_OPAD)
  );
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_BMUX = CLBLL_L_X2Y115_SLICE_X1Y115_B5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_CMUX = CLBLL_L_X2Y115_SLICE_X1Y115_C5Q;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_DMUX = CLBLL_L_X2Y115_SLICE_X1Y115_D5Q;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_AMUX = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BMUX = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_CMUX = CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_AMUX = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_BMUX = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_AMUX = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_BMUX = CLBLL_L_X2Y122_SLICE_X1Y122_B5Q;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B = CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_AMUX = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_BMUX = CLBLL_L_X4Y114_SLICE_X4Y114_B5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_AMUX = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CMUX = CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_DMUX = CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AMUX = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AMUX = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_AMUX = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_DMUX = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_AMUX = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_AMUX = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_BMUX = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CMUX = CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AMUX = CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CMUX = CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_DMUX = CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_BMUX = CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AMUX = CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_BMUX = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CMUX = CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_DMUX = CLBLL_L_X4Y120_SLICE_X5Y120_D5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_AMUX = CLBLL_L_X4Y121_SLICE_X5Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_BMUX = CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_DMUX = CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_AMUX = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_BMUX = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_AMUX = CLBLL_L_X4Y122_SLICE_X5Y122_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_CMUX = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A = CLBLL_L_X52Y113_SLICE_X78Y113_AO6;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B = CLBLL_L_X52Y113_SLICE_X78Y113_BO6;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C = CLBLL_L_X52Y113_SLICE_X78Y113_CO6;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D = CLBLL_L_X52Y113_SLICE_X78Y113_DO6;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A = CLBLL_L_X52Y113_SLICE_X79Y113_AO6;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B = CLBLL_L_X52Y113_SLICE_X79Y113_BO6;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C = CLBLL_L_X52Y113_SLICE_X79Y113_CO6;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D = CLBLL_L_X52Y113_SLICE_X79Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AMUX = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_BMUX = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AMUX = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_BMUX = CLBLM_R_X3Y113_SLICE_X3Y113_B5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_CMUX = CLBLM_R_X3Y113_SLICE_X3Y113_C5Q;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_DMUX = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AMUX = CLBLM_R_X3Y114_SLICE_X3Y114_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_BMUX = CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_CMUX = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AMUX = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_BMUX = CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CMUX = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_DMUX = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_AMUX = CLBLM_R_X3Y116_SLICE_X2Y116_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_BMUX = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_CMUX = CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_AMUX = CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_AMUX = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_BMUX = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_AMUX = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_AMUX = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_BMUX = CLBLM_R_X3Y119_SLICE_X3Y119_B5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AMUX = CLBLM_R_X3Y120_SLICE_X2Y120_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_CMUX = CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_DMUX = CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_BMUX = CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_CMUX = CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AMUX = CLBLM_R_X3Y121_SLICE_X2Y121_A5Q;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_BMUX = CLBLM_R_X3Y121_SLICE_X2Y121_B5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CMUX = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_DMUX = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AMUX = CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_BMUX = CLBLM_R_X3Y122_SLICE_X2Y122_B5Q;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_AMUX = CLBLM_R_X3Y122_SLICE_X3Y122_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_AMUX = CLBLM_R_X3Y123_SLICE_X2Y123_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AMUX = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_AMUX = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_BMUX = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_AMUX = CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_BMUX = CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_DMUX = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_BMUX = CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_AMUX = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_BMUX = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_DMUX = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_DMUX = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_DMUX = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_AMUX = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_BMUX = CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_AMUX = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_AMUX = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_AMUX = CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AMUX = CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_BMUX = CLBLM_R_X7Y120_SLICE_X8Y120_B5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CMUX = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_AMUX = CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CMUX = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_DMUX = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_O = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_O = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O = LIOB33_X0Y131_IOB_X0Y131_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_OQ = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_TQ = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_OQ = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_TQ = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_OQ = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_OQ = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_TQ = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_OQ = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_TQ = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_OQ = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_OQ = CLBLL_L_X52Y113_SLICE_X78Y113_AO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_TQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_OQ = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_OQ = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_OQ = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_OQ = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_OQ = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_TQ = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = 1'b1;
  assign RIOI3_X105Y109_OLOGIC_X1Y110_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_BX = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y109_OLOGIC_X1Y109_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = 1'b1;
  assign RIOB33_X105Y117_IOB_X1Y118_O = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign RIOB33_X105Y117_IOB_X1Y117_O = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AX = CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = CLBLL_L_X2Y120_SLICE_X1Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = 1'b1;
  assign RIOB33_X105Y119_IOB_X1Y119_O = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign RIOB33_X105Y119_IOB_X1Y120_O = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_B5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = CLBLM_R_X3Y119_SLICE_X3Y119_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AX = CLBLM_R_X3Y121_SLICE_X2Y121_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign RIOB33_X105Y121_IOB_X1Y121_O = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign RIOB33_X105Y121_IOB_X1Y122_O = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_BX = CLBLL_L_X2Y122_SLICE_X0Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLM_R_X3Y119_SLICE_X3Y119_B5Q;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLM_R_X3Y122_SLICE_X3Y122_A5Q;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_D1 = CLBLL_L_X52Y113_SLICE_X78Y113_AO6;
  assign RIOI3_X105Y111_OLOGIC_X1Y112_T1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_D1 = 1'b1;
  assign RIOI3_X105Y111_OLOGIC_X1Y111_T1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_AX = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AX = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_BX = 1'b0;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = CLBLM_R_X3Y121_SLICE_X2Y121_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = CLBLL_L_X4Y120_SLICE_X5Y120_D5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_B5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = CLBLL_L_X2Y122_SLICE_X0Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = CLBLM_R_X3Y122_SLICE_X2Y122_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = 1'b1;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_AX = CLBLM_R_X3Y123_SLICE_X2Y123_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLM_R_X3Y122_SLICE_X3Y122_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_AX = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_D = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_D = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = 1'b1;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_AX = CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AX = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_BX = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CX = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = CLBLL_L_X4Y120_SLICE_X5Y120_DQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_AX = CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = CLBLL_L_X2Y115_SLICE_X1Y115_B5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_D = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_D = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X7Y120_SLICE_X8Y120_B5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_R_X7Y120_SLICE_X8Y120_B5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_B5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_AX = CLBLM_R_X3Y120_SLICE_X2Y120_A5Q;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_BX = CLBLL_L_X2Y120_SLICE_X1Y120_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_AX = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_BX = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BX = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = CLBLL_L_X4Y114_SLICE_X4Y114_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_AX = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = CLBLM_R_X3Y121_SLICE_X2Y121_A5Q;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = CLBLL_L_X2Y122_SLICE_X0Y122_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = CLBLM_R_X3Y119_SLICE_X3Y119_B5Q;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = 1'b1;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_D = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = CLBLL_L_X4Y113_SLICE_X5Y113_DQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = 1'b1;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = CLBLL_L_X2Y122_SLICE_X0Y122_BQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_D5Q;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = CLBLM_R_X3Y122_SLICE_X2Y122_B5Q;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = CLBLL_L_X2Y122_SLICE_X1Y122_B5Q;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_BX = CLBLL_L_X2Y122_SLICE_X1Y122_CQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_CX = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = CLBLL_L_X4Y114_SLICE_X4Y114_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = CLBLL_L_X4Y114_SLICE_X4Y114_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = 1'b1;
  assign RIOI3_SING_X105Y100_OLOGIC_X1Y100_T1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_A6 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_B6 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_C6 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X78Y113_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_A6 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D1 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D2 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D3 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D4 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D5 = 1'b1;
  assign CLBLL_L_X52Y113_SLICE_X79Y113_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y108_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_D1 = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign RIOI3_TBYTESRC_X105Y107_OLOGIC_X1Y107_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLL_L_X2Y115_SLICE_X1Y115_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X3Y116_SLICE_X2Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_DQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLL_L_X4Y113_SLICE_X5Y113_DQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLL_L_X2Y115_SLICE_X1Y115_B5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AX = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_B5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CX = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_AX = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CX = CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_DX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = CLBLM_R_X3Y113_SLICE_X3Y113_CQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLM_R_X3Y113_SLICE_X3Y113_B5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLL_L_X2Y115_SLICE_X1Y115_D5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = CLBLL_L_X2Y115_SLICE_X1Y115_C5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLM_R_X3Y114_SLICE_X3Y114_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLM_R_X3Y113_SLICE_X3Y113_CQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = CLBLL_L_X2Y115_SLICE_X1Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = CLBLL_L_X2Y115_SLICE_X1Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = CLBLL_L_X2Y115_SLICE_X1Y115_C5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AX = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLM_R_X3Y114_SLICE_X3Y114_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLL_L_X2Y115_SLICE_X0Y115_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = CLBLM_R_X3Y113_SLICE_X3Y113_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = CLBLL_L_X2Y115_SLICE_X0Y115_CQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = CLBLL_L_X2Y115_SLICE_X0Y115_A5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A3 = CLBLM_R_X3Y122_SLICE_X2Y122_B5Q;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D2 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D3 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D4 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D5 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_AX = CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = CLBLM_R_X5Y121_SLICE_X6Y121_D5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_DQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_AX = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_AX = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y102_T1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = 1'b1;
  assign RIOI3_X105Y101_OLOGIC_X1Y101_T1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign RIOB33_X105Y101_IOB_X1Y101_O = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign RIOB33_X105Y101_IOB_X1Y102_O = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_AX = CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = CLBLM_R_X3Y120_SLICE_X2Y120_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = 1'b1;
  assign RIOB33_X105Y103_IOB_X1Y103_O = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign RIOB33_X105Y103_IOB_X1Y104_O = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AX = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_BX = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AX = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AX = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = CLBLL_L_X4Y114_SLICE_X5Y114_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOB33_X105Y105_IOB_X1Y106_O = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign RIOB33_X105Y105_IOB_X1Y105_O = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_BX = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLM_R_X3Y114_SLICE_X3Y114_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_CX = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLM_R_X3Y116_SLICE_X2Y116_DQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AX = CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign RIOI3_X105Y103_OLOGIC_X1Y104_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_D1 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign RIOI3_X105Y103_OLOGIC_X1Y103_T1 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLL_L_X4Y121_SLICE_X5Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_AX = CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOB33_X105Y107_IOB_X1Y108_O = 1'b1;
  assign RIOB33_X105Y107_IOB_X1Y107_O = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLL_L_X2Y115_SLICE_X1Y115_D5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AX = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = CLBLM_R_X3Y113_SLICE_X3Y113_C5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_BX = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLL_L_X2Y115_SLICE_X1Y115_DQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLM_R_X3Y113_SLICE_X3Y113_CQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AX = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = CLBLL_L_X2Y115_SLICE_X1Y115_C5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_BX = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CX = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLM_R_X3Y114_SLICE_X2Y114_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_AX = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = CLBLL_L_X4Y122_SLICE_X5Y122_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_CX = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_AX = CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_BX = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = CLBLL_L_X4Y122_SLICE_X4Y122_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = CLBLM_R_X5Y121_SLICE_X6Y121_CQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOB33_X105Y109_IOB_X1Y110_O = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign RIOB33_X105Y109_IOB_X1Y109_O = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = CLBLM_R_X3Y113_SLICE_X3Y113_C5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = CLBLL_L_X2Y115_SLICE_X1Y115_CQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_AX = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLL_L_X2Y115_SLICE_X1Y115_CQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_C5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = CLBLM_R_X3Y113_SLICE_X2Y113_CQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = CLBLM_R_X3Y113_SLICE_X3Y113_B5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = CLBLM_R_X3Y117_SLICE_X2Y117_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_DQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = CLBLL_L_X2Y115_SLICE_X0Y115_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign RIOI3_X105Y105_OLOGIC_X1Y106_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign RIOB33_X105Y111_IOB_X1Y112_O = CLBLL_L_X52Y113_SLICE_X78Y113_AO6;
  assign RIOB33_X105Y111_IOB_X1Y111_O = 1'b1;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign RIOI3_X105Y105_OLOGIC_X1Y105_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y114_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  assign RIOI3_TBYTETERM_X105Y113_OLOGIC_X1Y113_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = CLBLL_L_X4Y114_SLICE_X5Y114_BQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = CLBLL_L_X2Y115_SLICE_X1Y115_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = CLBLM_R_X3Y119_SLICE_X3Y119_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = CLBLL_L_X2Y115_SLICE_X1Y115_D5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = CLBLL_L_X2Y115_SLICE_X0Y115_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = 1'b1;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = CLBLM_R_X3Y116_SLICE_X2Y116_DQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_SR = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOB33_X105Y113_IOB_X1Y114_O = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign RIOB33_X105Y113_IOB_X1Y113_O = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_A5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_B5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = 1'b1;
  assign RIOB33_SING_X105Y100_IOB_X1Y100_O = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = 1'b1;
  assign RIOB33_X105Y115_IOB_X1Y116_O = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign RIOB33_X105Y115_IOB_X1Y115_O = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
endmodule
